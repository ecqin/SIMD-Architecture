//===================================================================
// Filename: harmonica_tracker_pred.sv
// Author: Eric Qin
// Purpose: Verification Module (test debugger)
//===================================================================


// Under Development
// TODO List
// 1) MACRO to get essential values in a readable form (non-synthesizable) // TODO
// 2) Print out of the register files based on thre warp and thread ID to read
// 3) Also serves as a checker and print out potential failed cases and timestamp
// 4) Look into tasks and interfaces
// 5) Make it generic to the point that timing changes doesnt affect the output as much
// FIXME -> code structure not efficient, too lengthy


`include "harmonica_cfg.sv" 

module harmonica_tracker_pred(
  input logic clk,
  // FIXME --> very wordy, not efficient
  // Interfaces? tasks? structs? need to look into this in the future
/*
  generate
    genvar GPR_index;
    for (GPR_index=0; GPR_index<NUM_TOTAL_THREADS; GPR_index=GPR_index+1) begin
      input logic [63:0] .NAME("GPR" + GPR_index)  [0:31];
    end
  endgenerate
*/
  input logic [63:0] PRED0 [0:31],
  input logic [63:0] PRED1 [0:31],
  input logic [63:0] PRED2 [0:31],
  input logic [63:0] PRED3 [0:31],
  input logic [63:0] PRED4 [0:31],
  input logic [63:0] PRED5 [0:31],
  input logic [63:0] PRED6 [0:31],
  input logic [63:0] PRED7 [0:31],
  input logic [63:0] PRED8 [0:31],
  input logic [63:0] PRED9 [0:31],
  input logic [63:0] PRED10 [0:31],
  input logic [63:0] PRED11 [0:31],
  input logic [63:0] PRED12 [0:31],
  input logic [63:0] PRED13 [0:31],
  input logic [63:0] PRED14 [0:31],
  input logic [63:0] PRED15 [0:31],
  input logic [63:0] PRED16 [0:31],
  input logic [63:0] PRED17 [0:31],
  input logic [63:0] PRED18 [0:31],
  input logic [63:0] PRED19 [0:31],
  input logic [63:0] PRED20 [0:31],
  input logic [63:0] PRED21 [0:31],
  input logic [63:0] PRED22 [0:31],
  input logic [63:0] PRED23 [0:31],
  input logic [63:0] PRED24 [0:31],
  input logic [63:0] PRED25 [0:31],
  input logic [63:0] PRED26 [0:31],
  input logic [63:0] PRED27 [0:31],
  input logic [63:0] PRED28 [0:31],
  input logic [63:0] PRED29 [0:31],
  input logic [63:0] PRED30 [0:31],
  input logic [63:0] PRED31 [0:31],
  input logic [63:0] PRED32 [0:31],
  input logic [63:0] PRED33 [0:31],
  input logic [63:0] PRED34 [0:31],
  input logic [63:0] PRED35 [0:31],
  input logic [63:0] PRED36 [0:31],
  input logic [63:0] PRED37 [0:31],
  input logic [63:0] PRED38 [0:31],
  input logic [63:0] PRED39 [0:31],
  input logic [63:0] PRED40 [0:31],
  input logic [63:0] PRED41 [0:31],
  input logic [63:0] PRED42 [0:31],
  input logic [63:0] PRED43 [0:31],
  input logic [63:0] PRED44 [0:31],
  input logic [63:0] PRED45 [0:31],
  input logic [63:0] PRED46 [0:31],
  input logic [63:0] PRED47 [0:31],
  input logic [63:0] PRED48 [0:31],
  input logic [63:0] PRED49 [0:31],
  input logic [63:0] PRED50 [0:31],
  input logic [63:0] PRED51 [0:31],
  input logic [63:0] PRED52 [0:31],
  input logic [63:0] PRED53 [0:31],
  input logic [63:0] PRED54 [0:31],
  input logic [63:0] PRED55 [0:31],
  input logic [63:0] PRED56 [0:31],
  input logic [63:0] PRED57 [0:31],
  input logic [63:0] PRED58 [0:31],
  input logic [63:0] PRED59 [0:31],
  input logic [63:0] PRED60 [0:31],
  input logic [63:0] PRED61 [0:31],
  input logic [63:0] PRED62 [0:31],
  input logic [63:0] PRED63 [0:31]
);

  integer f, i;
  // Initialize 2-entry buffers for comparison....

  // All register entry in all register files, code bloat. FIXME please, must be a better way, genvar???? 
  // 64 * 32 lol........
  logic [63:0] PRED0_0_buffer [0:1];
  logic [63:0] PRED0_1_buffer [0:1];
  logic [63:0] PRED0_2_buffer [0:1];
  logic [63:0] PRED0_3_buffer [0:1];
  logic [63:0] PRED0_4_buffer [0:1];
  logic [63:0] PRED0_5_buffer [0:1];
  logic [63:0] PRED0_6_buffer [0:1];
  logic [63:0] PRED0_7_buffer [0:1];
  logic [63:0] PRED0_8_buffer [0:1];
  logic [63:0] PRED0_9_buffer [0:1];
  logic [63:0] PRED0_10_buffer [0:1];
  logic [63:0] PRED0_11_buffer [0:1];
  logic [63:0] PRED0_12_buffer [0:1];
  logic [63:0] PRED0_13_buffer [0:1];
  logic [63:0] PRED0_14_buffer [0:1];
  logic [63:0] PRED0_15_buffer [0:1];
  logic [63:0] PRED0_16_buffer [0:1];
  logic [63:0] PRED0_17_buffer [0:1];
  logic [63:0] PRED0_18_buffer [0:1];
  logic [63:0] PRED0_19_buffer [0:1];
  logic [63:0] PRED0_20_buffer [0:1];
  logic [63:0] PRED0_21_buffer [0:1];
  logic [63:0] PRED0_22_buffer [0:1];
  logic [63:0] PRED0_23_buffer [0:1];
  logic [63:0] PRED0_24_buffer [0:1];
  logic [63:0] PRED0_25_buffer [0:1];
  logic [63:0] PRED0_26_buffer [0:1];
  logic [63:0] PRED0_27_buffer [0:1];
  logic [63:0] PRED0_28_buffer [0:1];
  logic [63:0] PRED0_29_buffer [0:1];
  logic [63:0] PRED0_30_buffer [0:1];
  logic [63:0] PRED0_31_buffer [0:1];
  logic [63:0] PRED1_0_buffer [0:1];
  logic [63:0] PRED1_1_buffer [0:1];
  logic [63:0] PRED1_2_buffer [0:1];
  logic [63:0] PRED1_3_buffer [0:1];
  logic [63:0] PRED1_4_buffer [0:1];
  logic [63:0] PRED1_5_buffer [0:1];
  logic [63:0] PRED1_6_buffer [0:1];
  logic [63:0] PRED1_7_buffer [0:1];
  logic [63:0] PRED1_8_buffer [0:1];
  logic [63:0] PRED1_9_buffer [0:1];
  logic [63:0] PRED1_10_buffer [0:1];
  logic [63:0] PRED1_11_buffer [0:1];
  logic [63:0] PRED1_12_buffer [0:1];
  logic [63:0] PRED1_13_buffer [0:1];
  logic [63:0] PRED1_14_buffer [0:1];
  logic [63:0] PRED1_15_buffer [0:1];
  logic [63:0] PRED1_16_buffer [0:1];
  logic [63:0] PRED1_17_buffer [0:1];
  logic [63:0] PRED1_18_buffer [0:1];
  logic [63:0] PRED1_19_buffer [0:1];
  logic [63:0] PRED1_20_buffer [0:1];
  logic [63:0] PRED1_21_buffer [0:1];
  logic [63:0] PRED1_22_buffer [0:1];
  logic [63:0] PRED1_23_buffer [0:1];
  logic [63:0] PRED1_24_buffer [0:1];
  logic [63:0] PRED1_25_buffer [0:1];
  logic [63:0] PRED1_26_buffer [0:1];
  logic [63:0] PRED1_27_buffer [0:1];
  logic [63:0] PRED1_28_buffer [0:1];
  logic [63:0] PRED1_29_buffer [0:1];
  logic [63:0] PRED1_30_buffer [0:1];
  logic [63:0] PRED1_31_buffer [0:1];
  logic [63:0] PRED2_0_buffer [0:1];
  logic [63:0] PRED2_1_buffer [0:1];
  logic [63:0] PRED2_2_buffer [0:1];
  logic [63:0] PRED2_3_buffer [0:1];
  logic [63:0] PRED2_4_buffer [0:1];
  logic [63:0] PRED2_5_buffer [0:1];
  logic [63:0] PRED2_6_buffer [0:1];
  logic [63:0] PRED2_7_buffer [0:1];
  logic [63:0] PRED2_8_buffer [0:1];
  logic [63:0] PRED2_9_buffer [0:1];
  logic [63:0] PRED2_10_buffer [0:1];
  logic [63:0] PRED2_11_buffer [0:1];
  logic [63:0] PRED2_12_buffer [0:1];
  logic [63:0] PRED2_13_buffer [0:1];
  logic [63:0] PRED2_14_buffer [0:1];
  logic [63:0] PRED2_15_buffer [0:1];
  logic [63:0] PRED2_16_buffer [0:1];
  logic [63:0] PRED2_17_buffer [0:1];
  logic [63:0] PRED2_18_buffer [0:1];
  logic [63:0] PRED2_19_buffer [0:1];
  logic [63:0] PRED2_20_buffer [0:1];
  logic [63:0] PRED2_21_buffer [0:1];
  logic [63:0] PRED2_22_buffer [0:1];
  logic [63:0] PRED2_23_buffer [0:1];
  logic [63:0] PRED2_24_buffer [0:1];
  logic [63:0] PRED2_25_buffer [0:1];
  logic [63:0] PRED2_26_buffer [0:1];
  logic [63:0] PRED2_27_buffer [0:1];
  logic [63:0] PRED2_28_buffer [0:1];
  logic [63:0] PRED2_29_buffer [0:1];
  logic [63:0] PRED2_30_buffer [0:1];
  logic [63:0] PRED2_31_buffer [0:1];
  logic [63:0] PRED3_0_buffer [0:1];
  logic [63:0] PRED3_1_buffer [0:1];
  logic [63:0] PRED3_2_buffer [0:1];
  logic [63:0] PRED3_3_buffer [0:1];
  logic [63:0] PRED3_4_buffer [0:1];
  logic [63:0] PRED3_5_buffer [0:1];
  logic [63:0] PRED3_6_buffer [0:1];
  logic [63:0] PRED3_7_buffer [0:1];
  logic [63:0] PRED3_8_buffer [0:1];
  logic [63:0] PRED3_9_buffer [0:1];
  logic [63:0] PRED3_10_buffer [0:1];
  logic [63:0] PRED3_11_buffer [0:1];
  logic [63:0] PRED3_12_buffer [0:1];
  logic [63:0] PRED3_13_buffer [0:1];
  logic [63:0] PRED3_14_buffer [0:1];
  logic [63:0] PRED3_15_buffer [0:1];
  logic [63:0] PRED3_16_buffer [0:1];
  logic [63:0] PRED3_17_buffer [0:1];
  logic [63:0] PRED3_18_buffer [0:1];
  logic [63:0] PRED3_19_buffer [0:1];
  logic [63:0] PRED3_20_buffer [0:1];
  logic [63:0] PRED3_21_buffer [0:1];
  logic [63:0] PRED3_22_buffer [0:1];
  logic [63:0] PRED3_23_buffer [0:1];
  logic [63:0] PRED3_24_buffer [0:1];
  logic [63:0] PRED3_25_buffer [0:1];
  logic [63:0] PRED3_26_buffer [0:1];
  logic [63:0] PRED3_27_buffer [0:1];
  logic [63:0] PRED3_28_buffer [0:1];
  logic [63:0] PRED3_29_buffer [0:1];
  logic [63:0] PRED3_30_buffer [0:1];
  logic [63:0] PRED3_31_buffer [0:1];
  logic [63:0] PRED4_0_buffer [0:1];
  logic [63:0] PRED4_1_buffer [0:1];
  logic [63:0] PRED4_2_buffer [0:1];
  logic [63:0] PRED4_3_buffer [0:1];
  logic [63:0] PRED4_4_buffer [0:1];
  logic [63:0] PRED4_5_buffer [0:1];
  logic [63:0] PRED4_6_buffer [0:1];
  logic [63:0] PRED4_7_buffer [0:1];
  logic [63:0] PRED4_8_buffer [0:1];
  logic [63:0] PRED4_9_buffer [0:1];
  logic [63:0] PRED4_10_buffer [0:1];
  logic [63:0] PRED4_11_buffer [0:1];
  logic [63:0] PRED4_12_buffer [0:1];
  logic [63:0] PRED4_13_buffer [0:1];
  logic [63:0] PRED4_14_buffer [0:1];
  logic [63:0] PRED4_15_buffer [0:1];
  logic [63:0] PRED4_16_buffer [0:1];
  logic [63:0] PRED4_17_buffer [0:1];
  logic [63:0] PRED4_18_buffer [0:1];
  logic [63:0] PRED4_19_buffer [0:1];
  logic [63:0] PRED4_20_buffer [0:1];
  logic [63:0] PRED4_21_buffer [0:1];
  logic [63:0] PRED4_22_buffer [0:1];
  logic [63:0] PRED4_23_buffer [0:1];
  logic [63:0] PRED4_24_buffer [0:1];
  logic [63:0] PRED4_25_buffer [0:1];
  logic [63:0] PRED4_26_buffer [0:1];
  logic [63:0] PRED4_27_buffer [0:1];
  logic [63:0] PRED4_28_buffer [0:1];
  logic [63:0] PRED4_29_buffer [0:1];
  logic [63:0] PRED4_30_buffer [0:1];
  logic [63:0] PRED4_31_buffer [0:1];
  logic [63:0] PRED5_0_buffer [0:1];
  logic [63:0] PRED5_1_buffer [0:1];
  logic [63:0] PRED5_2_buffer [0:1];
  logic [63:0] PRED5_3_buffer [0:1];
  logic [63:0] PRED5_4_buffer [0:1];
  logic [63:0] PRED5_5_buffer [0:1];
  logic [63:0] PRED5_6_buffer [0:1];
  logic [63:0] PRED5_7_buffer [0:1];
  logic [63:0] PRED5_8_buffer [0:1];
  logic [63:0] PRED5_9_buffer [0:1];
  logic [63:0] PRED5_10_buffer [0:1];
  logic [63:0] PRED5_11_buffer [0:1];
  logic [63:0] PRED5_12_buffer [0:1];
  logic [63:0] PRED5_13_buffer [0:1];
  logic [63:0] PRED5_14_buffer [0:1];
  logic [63:0] PRED5_15_buffer [0:1];
  logic [63:0] PRED5_16_buffer [0:1];
  logic [63:0] PRED5_17_buffer [0:1];
  logic [63:0] PRED5_18_buffer [0:1];
  logic [63:0] PRED5_19_buffer [0:1];
  logic [63:0] PRED5_20_buffer [0:1];
  logic [63:0] PRED5_21_buffer [0:1];
  logic [63:0] PRED5_22_buffer [0:1];
  logic [63:0] PRED5_23_buffer [0:1];
  logic [63:0] PRED5_24_buffer [0:1];
  logic [63:0] PRED5_25_buffer [0:1];
  logic [63:0] PRED5_26_buffer [0:1];
  logic [63:0] PRED5_27_buffer [0:1];
  logic [63:0] PRED5_28_buffer [0:1];
  logic [63:0] PRED5_29_buffer [0:1];
  logic [63:0] PRED5_30_buffer [0:1];
  logic [63:0] PRED5_31_buffer [0:1];
  logic [63:0] PRED6_0_buffer [0:1];
  logic [63:0] PRED6_1_buffer [0:1];
  logic [63:0] PRED6_2_buffer [0:1];
  logic [63:0] PRED6_3_buffer [0:1];
  logic [63:0] PRED6_4_buffer [0:1];
  logic [63:0] PRED6_5_buffer [0:1];
  logic [63:0] PRED6_6_buffer [0:1];
  logic [63:0] PRED6_7_buffer [0:1];
  logic [63:0] PRED6_8_buffer [0:1];
  logic [63:0] PRED6_9_buffer [0:1];
  logic [63:0] PRED6_10_buffer [0:1];
  logic [63:0] PRED6_11_buffer [0:1];
  logic [63:0] PRED6_12_buffer [0:1];
  logic [63:0] PRED6_13_buffer [0:1];
  logic [63:0] PRED6_14_buffer [0:1];
  logic [63:0] PRED6_15_buffer [0:1];
  logic [63:0] PRED6_16_buffer [0:1];
  logic [63:0] PRED6_17_buffer [0:1];
  logic [63:0] PRED6_18_buffer [0:1];
  logic [63:0] PRED6_19_buffer [0:1];
  logic [63:0] PRED6_20_buffer [0:1];
  logic [63:0] PRED6_21_buffer [0:1];
  logic [63:0] PRED6_22_buffer [0:1];
  logic [63:0] PRED6_23_buffer [0:1];
  logic [63:0] PRED6_24_buffer [0:1];
  logic [63:0] PRED6_25_buffer [0:1];
  logic [63:0] PRED6_26_buffer [0:1];
  logic [63:0] PRED6_27_buffer [0:1];
  logic [63:0] PRED6_28_buffer [0:1];
  logic [63:0] PRED6_29_buffer [0:1];
  logic [63:0] PRED6_30_buffer [0:1];
  logic [63:0] PRED6_31_buffer [0:1];
  logic [63:0] PRED7_0_buffer [0:1];
  logic [63:0] PRED7_1_buffer [0:1];
  logic [63:0] PRED7_2_buffer [0:1];
  logic [63:0] PRED7_3_buffer [0:1];
  logic [63:0] PRED7_4_buffer [0:1];
  logic [63:0] PRED7_5_buffer [0:1];
  logic [63:0] PRED7_6_buffer [0:1];
  logic [63:0] PRED7_7_buffer [0:1];
  logic [63:0] PRED7_8_buffer [0:1];
  logic [63:0] PRED7_9_buffer [0:1];
  logic [63:0] PRED7_10_buffer [0:1];
  logic [63:0] PRED7_11_buffer [0:1];
  logic [63:0] PRED7_12_buffer [0:1];
  logic [63:0] PRED7_13_buffer [0:1];
  logic [63:0] PRED7_14_buffer [0:1];
  logic [63:0] PRED7_15_buffer [0:1];
  logic [63:0] PRED7_16_buffer [0:1];
  logic [63:0] PRED7_17_buffer [0:1];
  logic [63:0] PRED7_18_buffer [0:1];
  logic [63:0] PRED7_19_buffer [0:1];
  logic [63:0] PRED7_20_buffer [0:1];
  logic [63:0] PRED7_21_buffer [0:1];
  logic [63:0] PRED7_22_buffer [0:1];
  logic [63:0] PRED7_23_buffer [0:1];
  logic [63:0] PRED7_24_buffer [0:1];
  logic [63:0] PRED7_25_buffer [0:1];
  logic [63:0] PRED7_26_buffer [0:1];
  logic [63:0] PRED7_27_buffer [0:1];
  logic [63:0] PRED7_28_buffer [0:1];
  logic [63:0] PRED7_29_buffer [0:1];
  logic [63:0] PRED7_30_buffer [0:1];
  logic [63:0] PRED7_31_buffer [0:1];
  logic [63:0] PRED8_0_buffer [0:1];
  logic [63:0] PRED8_1_buffer [0:1];
  logic [63:0] PRED8_2_buffer [0:1];
  logic [63:0] PRED8_3_buffer [0:1];
  logic [63:0] PRED8_4_buffer [0:1];
  logic [63:0] PRED8_5_buffer [0:1];
  logic [63:0] PRED8_6_buffer [0:1];
  logic [63:0] PRED8_7_buffer [0:1];
  logic [63:0] PRED8_8_buffer [0:1];
  logic [63:0] PRED8_9_buffer [0:1];
  logic [63:0] PRED8_10_buffer [0:1];
  logic [63:0] PRED8_11_buffer [0:1];
  logic [63:0] PRED8_12_buffer [0:1];
  logic [63:0] PRED8_13_buffer [0:1];
  logic [63:0] PRED8_14_buffer [0:1];
  logic [63:0] PRED8_15_buffer [0:1];
  logic [63:0] PRED8_16_buffer [0:1];
  logic [63:0] PRED8_17_buffer [0:1];
  logic [63:0] PRED8_18_buffer [0:1];
  logic [63:0] PRED8_19_buffer [0:1];
  logic [63:0] PRED8_20_buffer [0:1];
  logic [63:0] PRED8_21_buffer [0:1];
  logic [63:0] PRED8_22_buffer [0:1];
  logic [63:0] PRED8_23_buffer [0:1];
  logic [63:0] PRED8_24_buffer [0:1];
  logic [63:0] PRED8_25_buffer [0:1];
  logic [63:0] PRED8_26_buffer [0:1];
  logic [63:0] PRED8_27_buffer [0:1];
  logic [63:0] PRED8_28_buffer [0:1];
  logic [63:0] PRED8_29_buffer [0:1];
  logic [63:0] PRED8_30_buffer [0:1];
  logic [63:0] PRED8_31_buffer [0:1];
  logic [63:0] PRED9_0_buffer [0:1];
  logic [63:0] PRED9_1_buffer [0:1];
  logic [63:0] PRED9_2_buffer [0:1];
  logic [63:0] PRED9_3_buffer [0:1];
  logic [63:0] PRED9_4_buffer [0:1];
  logic [63:0] PRED9_5_buffer [0:1];
  logic [63:0] PRED9_6_buffer [0:1];
  logic [63:0] PRED9_7_buffer [0:1];
  logic [63:0] PRED9_8_buffer [0:1];
  logic [63:0] PRED9_9_buffer [0:1];
  logic [63:0] PRED9_10_buffer [0:1];
  logic [63:0] PRED9_11_buffer [0:1];
  logic [63:0] PRED9_12_buffer [0:1];
  logic [63:0] PRED9_13_buffer [0:1];
  logic [63:0] PRED9_14_buffer [0:1];
  logic [63:0] PRED9_15_buffer [0:1];
  logic [63:0] PRED9_16_buffer [0:1];
  logic [63:0] PRED9_17_buffer [0:1];
  logic [63:0] PRED9_18_buffer [0:1];
  logic [63:0] PRED9_19_buffer [0:1];
  logic [63:0] PRED9_20_buffer [0:1];
  logic [63:0] PRED9_21_buffer [0:1];
  logic [63:0] PRED9_22_buffer [0:1];
  logic [63:0] PRED9_23_buffer [0:1];
  logic [63:0] PRED9_24_buffer [0:1];
  logic [63:0] PRED9_25_buffer [0:1];
  logic [63:0] PRED9_26_buffer [0:1];
  logic [63:0] PRED9_27_buffer [0:1];
  logic [63:0] PRED9_28_buffer [0:1];
  logic [63:0] PRED9_29_buffer [0:1];
  logic [63:0] PRED9_30_buffer [0:1];
  logic [63:0] PRED9_31_buffer [0:1];
  logic [63:0] PRED10_0_buffer [0:1];
  logic [63:0] PRED10_1_buffer [0:1];
  logic [63:0] PRED10_2_buffer [0:1];
  logic [63:0] PRED10_3_buffer [0:1];
  logic [63:0] PRED10_4_buffer [0:1];
  logic [63:0] PRED10_5_buffer [0:1];
  logic [63:0] PRED10_6_buffer [0:1];
  logic [63:0] PRED10_7_buffer [0:1];
  logic [63:0] PRED10_8_buffer [0:1];
  logic [63:0] PRED10_9_buffer [0:1];
  logic [63:0] PRED10_10_buffer [0:1];
  logic [63:0] PRED10_11_buffer [0:1];
  logic [63:0] PRED10_12_buffer [0:1];
  logic [63:0] PRED10_13_buffer [0:1];
  logic [63:0] PRED10_14_buffer [0:1];
  logic [63:0] PRED10_15_buffer [0:1];
  logic [63:0] PRED10_16_buffer [0:1];
  logic [63:0] PRED10_17_buffer [0:1];
  logic [63:0] PRED10_18_buffer [0:1];
  logic [63:0] PRED10_19_buffer [0:1];
  logic [63:0] PRED10_20_buffer [0:1];
  logic [63:0] PRED10_21_buffer [0:1];
  logic [63:0] PRED10_22_buffer [0:1];
  logic [63:0] PRED10_23_buffer [0:1];
  logic [63:0] PRED10_24_buffer [0:1];
  logic [63:0] PRED10_25_buffer [0:1];
  logic [63:0] PRED10_26_buffer [0:1];
  logic [63:0] PRED10_27_buffer [0:1];
  logic [63:0] PRED10_28_buffer [0:1];
  logic [63:0] PRED10_29_buffer [0:1];
  logic [63:0] PRED10_30_buffer [0:1];
  logic [63:0] PRED10_31_buffer [0:1];
  logic [63:0] PRED11_0_buffer [0:1];
  logic [63:0] PRED11_1_buffer [0:1];
  logic [63:0] PRED11_2_buffer [0:1];
  logic [63:0] PRED11_3_buffer [0:1];
  logic [63:0] PRED11_4_buffer [0:1];
  logic [63:0] PRED11_5_buffer [0:1];
  logic [63:0] PRED11_6_buffer [0:1];
  logic [63:0] PRED11_7_buffer [0:1];
  logic [63:0] PRED11_8_buffer [0:1];
  logic [63:0] PRED11_9_buffer [0:1];
  logic [63:0] PRED11_10_buffer [0:1];
  logic [63:0] PRED11_11_buffer [0:1];
  logic [63:0] PRED11_12_buffer [0:1];
  logic [63:0] PRED11_13_buffer [0:1];
  logic [63:0] PRED11_14_buffer [0:1];
  logic [63:0] PRED11_15_buffer [0:1];
  logic [63:0] PRED11_16_buffer [0:1];
  logic [63:0] PRED11_17_buffer [0:1];
  logic [63:0] PRED11_18_buffer [0:1];
  logic [63:0] PRED11_19_buffer [0:1];
  logic [63:0] PRED11_20_buffer [0:1];
  logic [63:0] PRED11_21_buffer [0:1];
  logic [63:0] PRED11_22_buffer [0:1];
  logic [63:0] PRED11_23_buffer [0:1];
  logic [63:0] PRED11_24_buffer [0:1];
  logic [63:0] PRED11_25_buffer [0:1];
  logic [63:0] PRED11_26_buffer [0:1];
  logic [63:0] PRED11_27_buffer [0:1];
  logic [63:0] PRED11_28_buffer [0:1];
  logic [63:0] PRED11_29_buffer [0:1];
  logic [63:0] PRED11_30_buffer [0:1];
  logic [63:0] PRED11_31_buffer [0:1];
  logic [63:0] PRED12_0_buffer [0:1];
  logic [63:0] PRED12_1_buffer [0:1];
  logic [63:0] PRED12_2_buffer [0:1];
  logic [63:0] PRED12_3_buffer [0:1];
  logic [63:0] PRED12_4_buffer [0:1];
  logic [63:0] PRED12_5_buffer [0:1];
  logic [63:0] PRED12_6_buffer [0:1];
  logic [63:0] PRED12_7_buffer [0:1];
  logic [63:0] PRED12_8_buffer [0:1];
  logic [63:0] PRED12_9_buffer [0:1];
  logic [63:0] PRED12_10_buffer [0:1];
  logic [63:0] PRED12_11_buffer [0:1];
  logic [63:0] PRED12_12_buffer [0:1];
  logic [63:0] PRED12_13_buffer [0:1];
  logic [63:0] PRED12_14_buffer [0:1];
  logic [63:0] PRED12_15_buffer [0:1];
  logic [63:0] PRED12_16_buffer [0:1];
  logic [63:0] PRED12_17_buffer [0:1];
  logic [63:0] PRED12_18_buffer [0:1];
  logic [63:0] PRED12_19_buffer [0:1];
  logic [63:0] PRED12_20_buffer [0:1];
  logic [63:0] PRED12_21_buffer [0:1];
  logic [63:0] PRED12_22_buffer [0:1];
  logic [63:0] PRED12_23_buffer [0:1];
  logic [63:0] PRED12_24_buffer [0:1];
  logic [63:0] PRED12_25_buffer [0:1];
  logic [63:0] PRED12_26_buffer [0:1];
  logic [63:0] PRED12_27_buffer [0:1];
  logic [63:0] PRED12_28_buffer [0:1];
  logic [63:0] PRED12_29_buffer [0:1];
  logic [63:0] PRED12_30_buffer [0:1];
  logic [63:0] PRED12_31_buffer [0:1];
  logic [63:0] PRED13_0_buffer [0:1];
  logic [63:0] PRED13_1_buffer [0:1];
  logic [63:0] PRED13_2_buffer [0:1];
  logic [63:0] PRED13_3_buffer [0:1];
  logic [63:0] PRED13_4_buffer [0:1];
  logic [63:0] PRED13_5_buffer [0:1];
  logic [63:0] PRED13_6_buffer [0:1];
  logic [63:0] PRED13_7_buffer [0:1];
  logic [63:0] PRED13_8_buffer [0:1];
  logic [63:0] PRED13_9_buffer [0:1];
  logic [63:0] PRED13_10_buffer [0:1];
  logic [63:0] PRED13_11_buffer [0:1];
  logic [63:0] PRED13_12_buffer [0:1];
  logic [63:0] PRED13_13_buffer [0:1];
  logic [63:0] PRED13_14_buffer [0:1];
  logic [63:0] PRED13_15_buffer [0:1];
  logic [63:0] PRED13_16_buffer [0:1];
  logic [63:0] PRED13_17_buffer [0:1];
  logic [63:0] PRED13_18_buffer [0:1];
  logic [63:0] PRED13_19_buffer [0:1];
  logic [63:0] PRED13_20_buffer [0:1];
  logic [63:0] PRED13_21_buffer [0:1];
  logic [63:0] PRED13_22_buffer [0:1];
  logic [63:0] PRED13_23_buffer [0:1];
  logic [63:0] PRED13_24_buffer [0:1];
  logic [63:0] PRED13_25_buffer [0:1];
  logic [63:0] PRED13_26_buffer [0:1];
  logic [63:0] PRED13_27_buffer [0:1];
  logic [63:0] PRED13_28_buffer [0:1];
  logic [63:0] PRED13_29_buffer [0:1];
  logic [63:0] PRED13_30_buffer [0:1];
  logic [63:0] PRED13_31_buffer [0:1];
  logic [63:0] PRED14_0_buffer [0:1];
  logic [63:0] PRED14_1_buffer [0:1];
  logic [63:0] PRED14_2_buffer [0:1];
  logic [63:0] PRED14_3_buffer [0:1];
  logic [63:0] PRED14_4_buffer [0:1];
  logic [63:0] PRED14_5_buffer [0:1];
  logic [63:0] PRED14_6_buffer [0:1];
  logic [63:0] PRED14_7_buffer [0:1];
  logic [63:0] PRED14_8_buffer [0:1];
  logic [63:0] PRED14_9_buffer [0:1];
  logic [63:0] PRED14_10_buffer [0:1];
  logic [63:0] PRED14_11_buffer [0:1];
  logic [63:0] PRED14_12_buffer [0:1];
  logic [63:0] PRED14_13_buffer [0:1];
  logic [63:0] PRED14_14_buffer [0:1];
  logic [63:0] PRED14_15_buffer [0:1];
  logic [63:0] PRED14_16_buffer [0:1];
  logic [63:0] PRED14_17_buffer [0:1];
  logic [63:0] PRED14_18_buffer [0:1];
  logic [63:0] PRED14_19_buffer [0:1];
  logic [63:0] PRED14_20_buffer [0:1];
  logic [63:0] PRED14_21_buffer [0:1];
  logic [63:0] PRED14_22_buffer [0:1];
  logic [63:0] PRED14_23_buffer [0:1];
  logic [63:0] PRED14_24_buffer [0:1];
  logic [63:0] PRED14_25_buffer [0:1];
  logic [63:0] PRED14_26_buffer [0:1];
  logic [63:0] PRED14_27_buffer [0:1];
  logic [63:0] PRED14_28_buffer [0:1];
  logic [63:0] PRED14_29_buffer [0:1];
  logic [63:0] PRED14_30_buffer [0:1];
  logic [63:0] PRED14_31_buffer [0:1];
  logic [63:0] PRED15_0_buffer [0:1];
  logic [63:0] PRED15_1_buffer [0:1];
  logic [63:0] PRED15_2_buffer [0:1];
  logic [63:0] PRED15_3_buffer [0:1];
  logic [63:0] PRED15_4_buffer [0:1];
  logic [63:0] PRED15_5_buffer [0:1];
  logic [63:0] PRED15_6_buffer [0:1];
  logic [63:0] PRED15_7_buffer [0:1];
  logic [63:0] PRED15_8_buffer [0:1];
  logic [63:0] PRED15_9_buffer [0:1];
  logic [63:0] PRED15_10_buffer [0:1];
  logic [63:0] PRED15_11_buffer [0:1];
  logic [63:0] PRED15_12_buffer [0:1];
  logic [63:0] PRED15_13_buffer [0:1];
  logic [63:0] PRED15_14_buffer [0:1];
  logic [63:0] PRED15_15_buffer [0:1];
  logic [63:0] PRED15_16_buffer [0:1];
  logic [63:0] PRED15_17_buffer [0:1];
  logic [63:0] PRED15_18_buffer [0:1];
  logic [63:0] PRED15_19_buffer [0:1];
  logic [63:0] PRED15_20_buffer [0:1];
  logic [63:0] PRED15_21_buffer [0:1];
  logic [63:0] PRED15_22_buffer [0:1];
  logic [63:0] PRED15_23_buffer [0:1];
  logic [63:0] PRED15_24_buffer [0:1];
  logic [63:0] PRED15_25_buffer [0:1];
  logic [63:0] PRED15_26_buffer [0:1];
  logic [63:0] PRED15_27_buffer [0:1];
  logic [63:0] PRED15_28_buffer [0:1];
  logic [63:0] PRED15_29_buffer [0:1];
  logic [63:0] PRED15_30_buffer [0:1];
  logic [63:0] PRED15_31_buffer [0:1];
  logic [63:0] PRED16_0_buffer [0:1];
  logic [63:0] PRED16_1_buffer [0:1];
  logic [63:0] PRED16_2_buffer [0:1];
  logic [63:0] PRED16_3_buffer [0:1];
  logic [63:0] PRED16_4_buffer [0:1];
  logic [63:0] PRED16_5_buffer [0:1];
  logic [63:0] PRED16_6_buffer [0:1];
  logic [63:0] PRED16_7_buffer [0:1];
  logic [63:0] PRED16_8_buffer [0:1];
  logic [63:0] PRED16_9_buffer [0:1];
  logic [63:0] PRED16_10_buffer [0:1];
  logic [63:0] PRED16_11_buffer [0:1];
  logic [63:0] PRED16_12_buffer [0:1];
  logic [63:0] PRED16_13_buffer [0:1];
  logic [63:0] PRED16_14_buffer [0:1];
  logic [63:0] PRED16_15_buffer [0:1];
  logic [63:0] PRED16_16_buffer [0:1];
  logic [63:0] PRED16_17_buffer [0:1];
  logic [63:0] PRED16_18_buffer [0:1];
  logic [63:0] PRED16_19_buffer [0:1];
  logic [63:0] PRED16_20_buffer [0:1];
  logic [63:0] PRED16_21_buffer [0:1];
  logic [63:0] PRED16_22_buffer [0:1];
  logic [63:0] PRED16_23_buffer [0:1];
  logic [63:0] PRED16_24_buffer [0:1];
  logic [63:0] PRED16_25_buffer [0:1];
  logic [63:0] PRED16_26_buffer [0:1];
  logic [63:0] PRED16_27_buffer [0:1];
  logic [63:0] PRED16_28_buffer [0:1];
  logic [63:0] PRED16_29_buffer [0:1];
  logic [63:0] PRED16_30_buffer [0:1];
  logic [63:0] PRED16_31_buffer [0:1];
  logic [63:0] PRED17_0_buffer [0:1];
  logic [63:0] PRED17_1_buffer [0:1];
  logic [63:0] PRED17_2_buffer [0:1];
  logic [63:0] PRED17_3_buffer [0:1];
  logic [63:0] PRED17_4_buffer [0:1];
  logic [63:0] PRED17_5_buffer [0:1];
  logic [63:0] PRED17_6_buffer [0:1];
  logic [63:0] PRED17_7_buffer [0:1];
  logic [63:0] PRED17_8_buffer [0:1];
  logic [63:0] PRED17_9_buffer [0:1];
  logic [63:0] PRED17_10_buffer [0:1];
  logic [63:0] PRED17_11_buffer [0:1];
  logic [63:0] PRED17_12_buffer [0:1];
  logic [63:0] PRED17_13_buffer [0:1];
  logic [63:0] PRED17_14_buffer [0:1];
  logic [63:0] PRED17_15_buffer [0:1];
  logic [63:0] PRED17_16_buffer [0:1];
  logic [63:0] PRED17_17_buffer [0:1];
  logic [63:0] PRED17_18_buffer [0:1];
  logic [63:0] PRED17_19_buffer [0:1];
  logic [63:0] PRED17_20_buffer [0:1];
  logic [63:0] PRED17_21_buffer [0:1];
  logic [63:0] PRED17_22_buffer [0:1];
  logic [63:0] PRED17_23_buffer [0:1];
  logic [63:0] PRED17_24_buffer [0:1];
  logic [63:0] PRED17_25_buffer [0:1];
  logic [63:0] PRED17_26_buffer [0:1];
  logic [63:0] PRED17_27_buffer [0:1];
  logic [63:0] PRED17_28_buffer [0:1];
  logic [63:0] PRED17_29_buffer [0:1];
  logic [63:0] PRED17_30_buffer [0:1];
  logic [63:0] PRED17_31_buffer [0:1];
  logic [63:0] PRED18_0_buffer [0:1];
  logic [63:0] PRED18_1_buffer [0:1];
  logic [63:0] PRED18_2_buffer [0:1];
  logic [63:0] PRED18_3_buffer [0:1];
  logic [63:0] PRED18_4_buffer [0:1];
  logic [63:0] PRED18_5_buffer [0:1];
  logic [63:0] PRED18_6_buffer [0:1];
  logic [63:0] PRED18_7_buffer [0:1];
  logic [63:0] PRED18_8_buffer [0:1];
  logic [63:0] PRED18_9_buffer [0:1];
  logic [63:0] PRED18_10_buffer [0:1];
  logic [63:0] PRED18_11_buffer [0:1];
  logic [63:0] PRED18_12_buffer [0:1];
  logic [63:0] PRED18_13_buffer [0:1];
  logic [63:0] PRED18_14_buffer [0:1];
  logic [63:0] PRED18_15_buffer [0:1];
  logic [63:0] PRED18_16_buffer [0:1];
  logic [63:0] PRED18_17_buffer [0:1];
  logic [63:0] PRED18_18_buffer [0:1];
  logic [63:0] PRED18_19_buffer [0:1];
  logic [63:0] PRED18_20_buffer [0:1];
  logic [63:0] PRED18_21_buffer [0:1];
  logic [63:0] PRED18_22_buffer [0:1];
  logic [63:0] PRED18_23_buffer [0:1];
  logic [63:0] PRED18_24_buffer [0:1];
  logic [63:0] PRED18_25_buffer [0:1];
  logic [63:0] PRED18_26_buffer [0:1];
  logic [63:0] PRED18_27_buffer [0:1];
  logic [63:0] PRED18_28_buffer [0:1];
  logic [63:0] PRED18_29_buffer [0:1];
  logic [63:0] PRED18_30_buffer [0:1];
  logic [63:0] PRED18_31_buffer [0:1];
  logic [63:0] PRED19_0_buffer [0:1];
  logic [63:0] PRED19_1_buffer [0:1];
  logic [63:0] PRED19_2_buffer [0:1];
  logic [63:0] PRED19_3_buffer [0:1];
  logic [63:0] PRED19_4_buffer [0:1];
  logic [63:0] PRED19_5_buffer [0:1];
  logic [63:0] PRED19_6_buffer [0:1];
  logic [63:0] PRED19_7_buffer [0:1];
  logic [63:0] PRED19_8_buffer [0:1];
  logic [63:0] PRED19_9_buffer [0:1];
  logic [63:0] PRED19_10_buffer [0:1];
  logic [63:0] PRED19_11_buffer [0:1];
  logic [63:0] PRED19_12_buffer [0:1];
  logic [63:0] PRED19_13_buffer [0:1];
  logic [63:0] PRED19_14_buffer [0:1];
  logic [63:0] PRED19_15_buffer [0:1];
  logic [63:0] PRED19_16_buffer [0:1];
  logic [63:0] PRED19_17_buffer [0:1];
  logic [63:0] PRED19_18_buffer [0:1];
  logic [63:0] PRED19_19_buffer [0:1];
  logic [63:0] PRED19_20_buffer [0:1];
  logic [63:0] PRED19_21_buffer [0:1];
  logic [63:0] PRED19_22_buffer [0:1];
  logic [63:0] PRED19_23_buffer [0:1];
  logic [63:0] PRED19_24_buffer [0:1];
  logic [63:0] PRED19_25_buffer [0:1];
  logic [63:0] PRED19_26_buffer [0:1];
  logic [63:0] PRED19_27_buffer [0:1];
  logic [63:0] PRED19_28_buffer [0:1];
  logic [63:0] PRED19_29_buffer [0:1];
  logic [63:0] PRED19_30_buffer [0:1];
  logic [63:0] PRED19_31_buffer [0:1];
  logic [63:0] PRED20_0_buffer [0:1];
  logic [63:0] PRED20_1_buffer [0:1];
  logic [63:0] PRED20_2_buffer [0:1];
  logic [63:0] PRED20_3_buffer [0:1];
  logic [63:0] PRED20_4_buffer [0:1];
  logic [63:0] PRED20_5_buffer [0:1];
  logic [63:0] PRED20_6_buffer [0:1];
  logic [63:0] PRED20_7_buffer [0:1];
  logic [63:0] PRED20_8_buffer [0:1];
  logic [63:0] PRED20_9_buffer [0:1];
  logic [63:0] PRED20_10_buffer [0:1];
  logic [63:0] PRED20_11_buffer [0:1];
  logic [63:0] PRED20_12_buffer [0:1];
  logic [63:0] PRED20_13_buffer [0:1];
  logic [63:0] PRED20_14_buffer [0:1];
  logic [63:0] PRED20_15_buffer [0:1];
  logic [63:0] PRED20_16_buffer [0:1];
  logic [63:0] PRED20_17_buffer [0:1];
  logic [63:0] PRED20_18_buffer [0:1];
  logic [63:0] PRED20_19_buffer [0:1];
  logic [63:0] PRED20_20_buffer [0:1];
  logic [63:0] PRED20_21_buffer [0:1];
  logic [63:0] PRED20_22_buffer [0:1];
  logic [63:0] PRED20_23_buffer [0:1];
  logic [63:0] PRED20_24_buffer [0:1];
  logic [63:0] PRED20_25_buffer [0:1];
  logic [63:0] PRED20_26_buffer [0:1];
  logic [63:0] PRED20_27_buffer [0:1];
  logic [63:0] PRED20_28_buffer [0:1];
  logic [63:0] PRED20_29_buffer [0:1];
  logic [63:0] PRED20_30_buffer [0:1];
  logic [63:0] PRED20_31_buffer [0:1];
  logic [63:0] PRED21_0_buffer [0:1];
  logic [63:0] PRED21_1_buffer [0:1];
  logic [63:0] PRED21_2_buffer [0:1];
  logic [63:0] PRED21_3_buffer [0:1];
  logic [63:0] PRED21_4_buffer [0:1];
  logic [63:0] PRED21_5_buffer [0:1];
  logic [63:0] PRED21_6_buffer [0:1];
  logic [63:0] PRED21_7_buffer [0:1];
  logic [63:0] PRED21_8_buffer [0:1];
  logic [63:0] PRED21_9_buffer [0:1];
  logic [63:0] PRED21_10_buffer [0:1];
  logic [63:0] PRED21_11_buffer [0:1];
  logic [63:0] PRED21_12_buffer [0:1];
  logic [63:0] PRED21_13_buffer [0:1];
  logic [63:0] PRED21_14_buffer [0:1];
  logic [63:0] PRED21_15_buffer [0:1];
  logic [63:0] PRED21_16_buffer [0:1];
  logic [63:0] PRED21_17_buffer [0:1];
  logic [63:0] PRED21_18_buffer [0:1];
  logic [63:0] PRED21_19_buffer [0:1];
  logic [63:0] PRED21_20_buffer [0:1];
  logic [63:0] PRED21_21_buffer [0:1];
  logic [63:0] PRED21_22_buffer [0:1];
  logic [63:0] PRED21_23_buffer [0:1];
  logic [63:0] PRED21_24_buffer [0:1];
  logic [63:0] PRED21_25_buffer [0:1];
  logic [63:0] PRED21_26_buffer [0:1];
  logic [63:0] PRED21_27_buffer [0:1];
  logic [63:0] PRED21_28_buffer [0:1];
  logic [63:0] PRED21_29_buffer [0:1];
  logic [63:0] PRED21_30_buffer [0:1];
  logic [63:0] PRED21_31_buffer [0:1];
  logic [63:0] PRED22_0_buffer [0:1];
  logic [63:0] PRED22_1_buffer [0:1];
  logic [63:0] PRED22_2_buffer [0:1];
  logic [63:0] PRED22_3_buffer [0:1];
  logic [63:0] PRED22_4_buffer [0:1];
  logic [63:0] PRED22_5_buffer [0:1];
  logic [63:0] PRED22_6_buffer [0:1];
  logic [63:0] PRED22_7_buffer [0:1];
  logic [63:0] PRED22_8_buffer [0:1];
  logic [63:0] PRED22_9_buffer [0:1];
  logic [63:0] PRED22_10_buffer [0:1];
  logic [63:0] PRED22_11_buffer [0:1];
  logic [63:0] PRED22_12_buffer [0:1];
  logic [63:0] PRED22_13_buffer [0:1];
  logic [63:0] PRED22_14_buffer [0:1];
  logic [63:0] PRED22_15_buffer [0:1];
  logic [63:0] PRED22_16_buffer [0:1];
  logic [63:0] PRED22_17_buffer [0:1];
  logic [63:0] PRED22_18_buffer [0:1];
  logic [63:0] PRED22_19_buffer [0:1];
  logic [63:0] PRED22_20_buffer [0:1];
  logic [63:0] PRED22_21_buffer [0:1];
  logic [63:0] PRED22_22_buffer [0:1];
  logic [63:0] PRED22_23_buffer [0:1];
  logic [63:0] PRED22_24_buffer [0:1];
  logic [63:0] PRED22_25_buffer [0:1];
  logic [63:0] PRED22_26_buffer [0:1];
  logic [63:0] PRED22_27_buffer [0:1];
  logic [63:0] PRED22_28_buffer [0:1];
  logic [63:0] PRED22_29_buffer [0:1];
  logic [63:0] PRED22_30_buffer [0:1];
  logic [63:0] PRED22_31_buffer [0:1];
  logic [63:0] PRED23_0_buffer [0:1];
  logic [63:0] PRED23_1_buffer [0:1];
  logic [63:0] PRED23_2_buffer [0:1];
  logic [63:0] PRED23_3_buffer [0:1];
  logic [63:0] PRED23_4_buffer [0:1];
  logic [63:0] PRED23_5_buffer [0:1];
  logic [63:0] PRED23_6_buffer [0:1];
  logic [63:0] PRED23_7_buffer [0:1];
  logic [63:0] PRED23_8_buffer [0:1];
  logic [63:0] PRED23_9_buffer [0:1];
  logic [63:0] PRED23_10_buffer [0:1];
  logic [63:0] PRED23_11_buffer [0:1];
  logic [63:0] PRED23_12_buffer [0:1];
  logic [63:0] PRED23_13_buffer [0:1];
  logic [63:0] PRED23_14_buffer [0:1];
  logic [63:0] PRED23_15_buffer [0:1];
  logic [63:0] PRED23_16_buffer [0:1];
  logic [63:0] PRED23_17_buffer [0:1];
  logic [63:0] PRED23_18_buffer [0:1];
  logic [63:0] PRED23_19_buffer [0:1];
  logic [63:0] PRED23_20_buffer [0:1];
  logic [63:0] PRED23_21_buffer [0:1];
  logic [63:0] PRED23_22_buffer [0:1];
  logic [63:0] PRED23_23_buffer [0:1];
  logic [63:0] PRED23_24_buffer [0:1];
  logic [63:0] PRED23_25_buffer [0:1];
  logic [63:0] PRED23_26_buffer [0:1];
  logic [63:0] PRED23_27_buffer [0:1];
  logic [63:0] PRED23_28_buffer [0:1];
  logic [63:0] PRED23_29_buffer [0:1];
  logic [63:0] PRED23_30_buffer [0:1];
  logic [63:0] PRED23_31_buffer [0:1];
  logic [63:0] PRED24_0_buffer [0:1];
  logic [63:0] PRED24_1_buffer [0:1];
  logic [63:0] PRED24_2_buffer [0:1];
  logic [63:0] PRED24_3_buffer [0:1];
  logic [63:0] PRED24_4_buffer [0:1];
  logic [63:0] PRED24_5_buffer [0:1];
  logic [63:0] PRED24_6_buffer [0:1];
  logic [63:0] PRED24_7_buffer [0:1];
  logic [63:0] PRED24_8_buffer [0:1];
  logic [63:0] PRED24_9_buffer [0:1];
  logic [63:0] PRED24_10_buffer [0:1];
  logic [63:0] PRED24_11_buffer [0:1];
  logic [63:0] PRED24_12_buffer [0:1];
  logic [63:0] PRED24_13_buffer [0:1];
  logic [63:0] PRED24_14_buffer [0:1];
  logic [63:0] PRED24_15_buffer [0:1];
  logic [63:0] PRED24_16_buffer [0:1];
  logic [63:0] PRED24_17_buffer [0:1];
  logic [63:0] PRED24_18_buffer [0:1];
  logic [63:0] PRED24_19_buffer [0:1];
  logic [63:0] PRED24_20_buffer [0:1];
  logic [63:0] PRED24_21_buffer [0:1];
  logic [63:0] PRED24_22_buffer [0:1];
  logic [63:0] PRED24_23_buffer [0:1];
  logic [63:0] PRED24_24_buffer [0:1];
  logic [63:0] PRED24_25_buffer [0:1];
  logic [63:0] PRED24_26_buffer [0:1];
  logic [63:0] PRED24_27_buffer [0:1];
  logic [63:0] PRED24_28_buffer [0:1];
  logic [63:0] PRED24_29_buffer [0:1];
  logic [63:0] PRED24_30_buffer [0:1];
  logic [63:0] PRED24_31_buffer [0:1];
  logic [63:0] PRED25_0_buffer [0:1];
  logic [63:0] PRED25_1_buffer [0:1];
  logic [63:0] PRED25_2_buffer [0:1];
  logic [63:0] PRED25_3_buffer [0:1];
  logic [63:0] PRED25_4_buffer [0:1];
  logic [63:0] PRED25_5_buffer [0:1];
  logic [63:0] PRED25_6_buffer [0:1];
  logic [63:0] PRED25_7_buffer [0:1];
  logic [63:0] PRED25_8_buffer [0:1];
  logic [63:0] PRED25_9_buffer [0:1];
  logic [63:0] PRED25_10_buffer [0:1];
  logic [63:0] PRED25_11_buffer [0:1];
  logic [63:0] PRED25_12_buffer [0:1];
  logic [63:0] PRED25_13_buffer [0:1];
  logic [63:0] PRED25_14_buffer [0:1];
  logic [63:0] PRED25_15_buffer [0:1];
  logic [63:0] PRED25_16_buffer [0:1];
  logic [63:0] PRED25_17_buffer [0:1];
  logic [63:0] PRED25_18_buffer [0:1];
  logic [63:0] PRED25_19_buffer [0:1];
  logic [63:0] PRED25_20_buffer [0:1];
  logic [63:0] PRED25_21_buffer [0:1];
  logic [63:0] PRED25_22_buffer [0:1];
  logic [63:0] PRED25_23_buffer [0:1];
  logic [63:0] PRED25_24_buffer [0:1];
  logic [63:0] PRED25_25_buffer [0:1];
  logic [63:0] PRED25_26_buffer [0:1];
  logic [63:0] PRED25_27_buffer [0:1];
  logic [63:0] PRED25_28_buffer [0:1];
  logic [63:0] PRED25_29_buffer [0:1];
  logic [63:0] PRED25_30_buffer [0:1];
  logic [63:0] PRED25_31_buffer [0:1];
  logic [63:0] PRED26_0_buffer [0:1];
  logic [63:0] PRED26_1_buffer [0:1];
  logic [63:0] PRED26_2_buffer [0:1];
  logic [63:0] PRED26_3_buffer [0:1];
  logic [63:0] PRED26_4_buffer [0:1];
  logic [63:0] PRED26_5_buffer [0:1];
  logic [63:0] PRED26_6_buffer [0:1];
  logic [63:0] PRED26_7_buffer [0:1];
  logic [63:0] PRED26_8_buffer [0:1];
  logic [63:0] PRED26_9_buffer [0:1];
  logic [63:0] PRED26_10_buffer [0:1];
  logic [63:0] PRED26_11_buffer [0:1];
  logic [63:0] PRED26_12_buffer [0:1];
  logic [63:0] PRED26_13_buffer [0:1];
  logic [63:0] PRED26_14_buffer [0:1];
  logic [63:0] PRED26_15_buffer [0:1];
  logic [63:0] PRED26_16_buffer [0:1];
  logic [63:0] PRED26_17_buffer [0:1];
  logic [63:0] PRED26_18_buffer [0:1];
  logic [63:0] PRED26_19_buffer [0:1];
  logic [63:0] PRED26_20_buffer [0:1];
  logic [63:0] PRED26_21_buffer [0:1];
  logic [63:0] PRED26_22_buffer [0:1];
  logic [63:0] PRED26_23_buffer [0:1];
  logic [63:0] PRED26_24_buffer [0:1];
  logic [63:0] PRED26_25_buffer [0:1];
  logic [63:0] PRED26_26_buffer [0:1];
  logic [63:0] PRED26_27_buffer [0:1];
  logic [63:0] PRED26_28_buffer [0:1];
  logic [63:0] PRED26_29_buffer [0:1];
  logic [63:0] PRED26_30_buffer [0:1];
  logic [63:0] PRED26_31_buffer [0:1];
  logic [63:0] PRED27_0_buffer [0:1];
  logic [63:0] PRED27_1_buffer [0:1];
  logic [63:0] PRED27_2_buffer [0:1];
  logic [63:0] PRED27_3_buffer [0:1];
  logic [63:0] PRED27_4_buffer [0:1];
  logic [63:0] PRED27_5_buffer [0:1];
  logic [63:0] PRED27_6_buffer [0:1];
  logic [63:0] PRED27_7_buffer [0:1];
  logic [63:0] PRED27_8_buffer [0:1];
  logic [63:0] PRED27_9_buffer [0:1];
  logic [63:0] PRED27_10_buffer [0:1];
  logic [63:0] PRED27_11_buffer [0:1];
  logic [63:0] PRED27_12_buffer [0:1];
  logic [63:0] PRED27_13_buffer [0:1];
  logic [63:0] PRED27_14_buffer [0:1];
  logic [63:0] PRED27_15_buffer [0:1];
  logic [63:0] PRED27_16_buffer [0:1];
  logic [63:0] PRED27_17_buffer [0:1];
  logic [63:0] PRED27_18_buffer [0:1];
  logic [63:0] PRED27_19_buffer [0:1];
  logic [63:0] PRED27_20_buffer [0:1];
  logic [63:0] PRED27_21_buffer [0:1];
  logic [63:0] PRED27_22_buffer [0:1];
  logic [63:0] PRED27_23_buffer [0:1];
  logic [63:0] PRED27_24_buffer [0:1];
  logic [63:0] PRED27_25_buffer [0:1];
  logic [63:0] PRED27_26_buffer [0:1];
  logic [63:0] PRED27_27_buffer [0:1];
  logic [63:0] PRED27_28_buffer [0:1];
  logic [63:0] PRED27_29_buffer [0:1];
  logic [63:0] PRED27_30_buffer [0:1];
  logic [63:0] PRED27_31_buffer [0:1];
  logic [63:0] PRED28_0_buffer [0:1];
  logic [63:0] PRED28_1_buffer [0:1];
  logic [63:0] PRED28_2_buffer [0:1];
  logic [63:0] PRED28_3_buffer [0:1];
  logic [63:0] PRED28_4_buffer [0:1];
  logic [63:0] PRED28_5_buffer [0:1];
  logic [63:0] PRED28_6_buffer [0:1];
  logic [63:0] PRED28_7_buffer [0:1];
  logic [63:0] PRED28_8_buffer [0:1];
  logic [63:0] PRED28_9_buffer [0:1];
  logic [63:0] PRED28_10_buffer [0:1];
  logic [63:0] PRED28_11_buffer [0:1];
  logic [63:0] PRED28_12_buffer [0:1];
  logic [63:0] PRED28_13_buffer [0:1];
  logic [63:0] PRED28_14_buffer [0:1];
  logic [63:0] PRED28_15_buffer [0:1];
  logic [63:0] PRED28_16_buffer [0:1];
  logic [63:0] PRED28_17_buffer [0:1];
  logic [63:0] PRED28_18_buffer [0:1];
  logic [63:0] PRED28_19_buffer [0:1];
  logic [63:0] PRED28_20_buffer [0:1];
  logic [63:0] PRED28_21_buffer [0:1];
  logic [63:0] PRED28_22_buffer [0:1];
  logic [63:0] PRED28_23_buffer [0:1];
  logic [63:0] PRED28_24_buffer [0:1];
  logic [63:0] PRED28_25_buffer [0:1];
  logic [63:0] PRED28_26_buffer [0:1];
  logic [63:0] PRED28_27_buffer [0:1];
  logic [63:0] PRED28_28_buffer [0:1];
  logic [63:0] PRED28_29_buffer [0:1];
  logic [63:0] PRED28_30_buffer [0:1];
  logic [63:0] PRED28_31_buffer [0:1];
  logic [63:0] PRED29_0_buffer [0:1];
  logic [63:0] PRED29_1_buffer [0:1];
  logic [63:0] PRED29_2_buffer [0:1];
  logic [63:0] PRED29_3_buffer [0:1];
  logic [63:0] PRED29_4_buffer [0:1];
  logic [63:0] PRED29_5_buffer [0:1];
  logic [63:0] PRED29_6_buffer [0:1];
  logic [63:0] PRED29_7_buffer [0:1];
  logic [63:0] PRED29_8_buffer [0:1];
  logic [63:0] PRED29_9_buffer [0:1];
  logic [63:0] PRED29_10_buffer [0:1];
  logic [63:0] PRED29_11_buffer [0:1];
  logic [63:0] PRED29_12_buffer [0:1];
  logic [63:0] PRED29_13_buffer [0:1];
  logic [63:0] PRED29_14_buffer [0:1];
  logic [63:0] PRED29_15_buffer [0:1];
  logic [63:0] PRED29_16_buffer [0:1];
  logic [63:0] PRED29_17_buffer [0:1];
  logic [63:0] PRED29_18_buffer [0:1];
  logic [63:0] PRED29_19_buffer [0:1];
  logic [63:0] PRED29_20_buffer [0:1];
  logic [63:0] PRED29_21_buffer [0:1];
  logic [63:0] PRED29_22_buffer [0:1];
  logic [63:0] PRED29_23_buffer [0:1];
  logic [63:0] PRED29_24_buffer [0:1];
  logic [63:0] PRED29_25_buffer [0:1];
  logic [63:0] PRED29_26_buffer [0:1];
  logic [63:0] PRED29_27_buffer [0:1];
  logic [63:0] PRED29_28_buffer [0:1];
  logic [63:0] PRED29_29_buffer [0:1];
  logic [63:0] PRED29_30_buffer [0:1];
  logic [63:0] PRED29_31_buffer [0:1];
  logic [63:0] PRED30_0_buffer [0:1];
  logic [63:0] PRED30_1_buffer [0:1];
  logic [63:0] PRED30_2_buffer [0:1];
  logic [63:0] PRED30_3_buffer [0:1];
  logic [63:0] PRED30_4_buffer [0:1];
  logic [63:0] PRED30_5_buffer [0:1];
  logic [63:0] PRED30_6_buffer [0:1];
  logic [63:0] PRED30_7_buffer [0:1];
  logic [63:0] PRED30_8_buffer [0:1];
  logic [63:0] PRED30_9_buffer [0:1];
  logic [63:0] PRED30_10_buffer [0:1];
  logic [63:0] PRED30_11_buffer [0:1];
  logic [63:0] PRED30_12_buffer [0:1];
  logic [63:0] PRED30_13_buffer [0:1];
  logic [63:0] PRED30_14_buffer [0:1];
  logic [63:0] PRED30_15_buffer [0:1];
  logic [63:0] PRED30_16_buffer [0:1];
  logic [63:0] PRED30_17_buffer [0:1];
  logic [63:0] PRED30_18_buffer [0:1];
  logic [63:0] PRED30_19_buffer [0:1];
  logic [63:0] PRED30_20_buffer [0:1];
  logic [63:0] PRED30_21_buffer [0:1];
  logic [63:0] PRED30_22_buffer [0:1];
  logic [63:0] PRED30_23_buffer [0:1];
  logic [63:0] PRED30_24_buffer [0:1];
  logic [63:0] PRED30_25_buffer [0:1];
  logic [63:0] PRED30_26_buffer [0:1];
  logic [63:0] PRED30_27_buffer [0:1];
  logic [63:0] PRED30_28_buffer [0:1];
  logic [63:0] PRED30_29_buffer [0:1];
  logic [63:0] PRED30_30_buffer [0:1];
  logic [63:0] PRED30_31_buffer [0:1];
  logic [63:0] PRED31_0_buffer [0:1];
  logic [63:0] PRED31_1_buffer [0:1];
  logic [63:0] PRED31_2_buffer [0:1];
  logic [63:0] PRED31_3_buffer [0:1];
  logic [63:0] PRED31_4_buffer [0:1];
  logic [63:0] PRED31_5_buffer [0:1];
  logic [63:0] PRED31_6_buffer [0:1];
  logic [63:0] PRED31_7_buffer [0:1];
  logic [63:0] PRED31_8_buffer [0:1];
  logic [63:0] PRED31_9_buffer [0:1];
  logic [63:0] PRED31_10_buffer [0:1];
  logic [63:0] PRED31_11_buffer [0:1];
  logic [63:0] PRED31_12_buffer [0:1];
  logic [63:0] PRED31_13_buffer [0:1];
  logic [63:0] PRED31_14_buffer [0:1];
  logic [63:0] PRED31_15_buffer [0:1];
  logic [63:0] PRED31_16_buffer [0:1];
  logic [63:0] PRED31_17_buffer [0:1];
  logic [63:0] PRED31_18_buffer [0:1];
  logic [63:0] PRED31_19_buffer [0:1];
  logic [63:0] PRED31_20_buffer [0:1];
  logic [63:0] PRED31_21_buffer [0:1];
  logic [63:0] PRED31_22_buffer [0:1];
  logic [63:0] PRED31_23_buffer [0:1];
  logic [63:0] PRED31_24_buffer [0:1];
  logic [63:0] PRED31_25_buffer [0:1];
  logic [63:0] PRED31_26_buffer [0:1];
  logic [63:0] PRED31_27_buffer [0:1];
  logic [63:0] PRED31_28_buffer [0:1];
  logic [63:0] PRED31_29_buffer [0:1];
  logic [63:0] PRED31_30_buffer [0:1];
  logic [63:0] PRED31_31_buffer [0:1];
  logic [63:0] PRED32_0_buffer [0:1];
  logic [63:0] PRED32_1_buffer [0:1];
  logic [63:0] PRED32_2_buffer [0:1];
  logic [63:0] PRED32_3_buffer [0:1];
  logic [63:0] PRED32_4_buffer [0:1];
  logic [63:0] PRED32_5_buffer [0:1];
  logic [63:0] PRED32_6_buffer [0:1];
  logic [63:0] PRED32_7_buffer [0:1];
  logic [63:0] PRED32_8_buffer [0:1];
  logic [63:0] PRED32_9_buffer [0:1];
  logic [63:0] PRED32_10_buffer [0:1];
  logic [63:0] PRED32_11_buffer [0:1];
  logic [63:0] PRED32_12_buffer [0:1];
  logic [63:0] PRED32_13_buffer [0:1];
  logic [63:0] PRED32_14_buffer [0:1];
  logic [63:0] PRED32_15_buffer [0:1];
  logic [63:0] PRED32_16_buffer [0:1];
  logic [63:0] PRED32_17_buffer [0:1];
  logic [63:0] PRED32_18_buffer [0:1];
  logic [63:0] PRED32_19_buffer [0:1];
  logic [63:0] PRED32_20_buffer [0:1];
  logic [63:0] PRED32_21_buffer [0:1];
  logic [63:0] PRED32_22_buffer [0:1];
  logic [63:0] PRED32_23_buffer [0:1];
  logic [63:0] PRED32_24_buffer [0:1];
  logic [63:0] PRED32_25_buffer [0:1];
  logic [63:0] PRED32_26_buffer [0:1];
  logic [63:0] PRED32_27_buffer [0:1];
  logic [63:0] PRED32_28_buffer [0:1];
  logic [63:0] PRED32_29_buffer [0:1];
  logic [63:0] PRED32_30_buffer [0:1];
  logic [63:0] PRED32_31_buffer [0:1];
  logic [63:0] PRED33_0_buffer [0:1];
  logic [63:0] PRED33_1_buffer [0:1];
  logic [63:0] PRED33_2_buffer [0:1];
  logic [63:0] PRED33_3_buffer [0:1];
  logic [63:0] PRED33_4_buffer [0:1];
  logic [63:0] PRED33_5_buffer [0:1];
  logic [63:0] PRED33_6_buffer [0:1];
  logic [63:0] PRED33_7_buffer [0:1];
  logic [63:0] PRED33_8_buffer [0:1];
  logic [63:0] PRED33_9_buffer [0:1];
  logic [63:0] PRED33_10_buffer [0:1];
  logic [63:0] PRED33_11_buffer [0:1];
  logic [63:0] PRED33_12_buffer [0:1];
  logic [63:0] PRED33_13_buffer [0:1];
  logic [63:0] PRED33_14_buffer [0:1];
  logic [63:0] PRED33_15_buffer [0:1];
  logic [63:0] PRED33_16_buffer [0:1];
  logic [63:0] PRED33_17_buffer [0:1];
  logic [63:0] PRED33_18_buffer [0:1];
  logic [63:0] PRED33_19_buffer [0:1];
  logic [63:0] PRED33_20_buffer [0:1];
  logic [63:0] PRED33_21_buffer [0:1];
  logic [63:0] PRED33_22_buffer [0:1];
  logic [63:0] PRED33_23_buffer [0:1];
  logic [63:0] PRED33_24_buffer [0:1];
  logic [63:0] PRED33_25_buffer [0:1];
  logic [63:0] PRED33_26_buffer [0:1];
  logic [63:0] PRED33_27_buffer [0:1];
  logic [63:0] PRED33_28_buffer [0:1];
  logic [63:0] PRED33_29_buffer [0:1];
  logic [63:0] PRED33_30_buffer [0:1];
  logic [63:0] PRED33_31_buffer [0:1];
  logic [63:0] PRED34_0_buffer [0:1];
  logic [63:0] PRED34_1_buffer [0:1];
  logic [63:0] PRED34_2_buffer [0:1];
  logic [63:0] PRED34_3_buffer [0:1];
  logic [63:0] PRED34_4_buffer [0:1];
  logic [63:0] PRED34_5_buffer [0:1];
  logic [63:0] PRED34_6_buffer [0:1];
  logic [63:0] PRED34_7_buffer [0:1];
  logic [63:0] PRED34_8_buffer [0:1];
  logic [63:0] PRED34_9_buffer [0:1];
  logic [63:0] PRED34_10_buffer [0:1];
  logic [63:0] PRED34_11_buffer [0:1];
  logic [63:0] PRED34_12_buffer [0:1];
  logic [63:0] PRED34_13_buffer [0:1];
  logic [63:0] PRED34_14_buffer [0:1];
  logic [63:0] PRED34_15_buffer [0:1];
  logic [63:0] PRED34_16_buffer [0:1];
  logic [63:0] PRED34_17_buffer [0:1];
  logic [63:0] PRED34_18_buffer [0:1];
  logic [63:0] PRED34_19_buffer [0:1];
  logic [63:0] PRED34_20_buffer [0:1];
  logic [63:0] PRED34_21_buffer [0:1];
  logic [63:0] PRED34_22_buffer [0:1];
  logic [63:0] PRED34_23_buffer [0:1];
  logic [63:0] PRED34_24_buffer [0:1];
  logic [63:0] PRED34_25_buffer [0:1];
  logic [63:0] PRED34_26_buffer [0:1];
  logic [63:0] PRED34_27_buffer [0:1];
  logic [63:0] PRED34_28_buffer [0:1];
  logic [63:0] PRED34_29_buffer [0:1];
  logic [63:0] PRED34_30_buffer [0:1];
  logic [63:0] PRED34_31_buffer [0:1];
  logic [63:0] PRED35_0_buffer [0:1];
  logic [63:0] PRED35_1_buffer [0:1];
  logic [63:0] PRED35_2_buffer [0:1];
  logic [63:0] PRED35_3_buffer [0:1];
  logic [63:0] PRED35_4_buffer [0:1];
  logic [63:0] PRED35_5_buffer [0:1];
  logic [63:0] PRED35_6_buffer [0:1];
  logic [63:0] PRED35_7_buffer [0:1];
  logic [63:0] PRED35_8_buffer [0:1];
  logic [63:0] PRED35_9_buffer [0:1];
  logic [63:0] PRED35_10_buffer [0:1];
  logic [63:0] PRED35_11_buffer [0:1];
  logic [63:0] PRED35_12_buffer [0:1];
  logic [63:0] PRED35_13_buffer [0:1];
  logic [63:0] PRED35_14_buffer [0:1];
  logic [63:0] PRED35_15_buffer [0:1];
  logic [63:0] PRED35_16_buffer [0:1];
  logic [63:0] PRED35_17_buffer [0:1];
  logic [63:0] PRED35_18_buffer [0:1];
  logic [63:0] PRED35_19_buffer [0:1];
  logic [63:0] PRED35_20_buffer [0:1];
  logic [63:0] PRED35_21_buffer [0:1];
  logic [63:0] PRED35_22_buffer [0:1];
  logic [63:0] PRED35_23_buffer [0:1];
  logic [63:0] PRED35_24_buffer [0:1];
  logic [63:0] PRED35_25_buffer [0:1];
  logic [63:0] PRED35_26_buffer [0:1];
  logic [63:0] PRED35_27_buffer [0:1];
  logic [63:0] PRED35_28_buffer [0:1];
  logic [63:0] PRED35_29_buffer [0:1];
  logic [63:0] PRED35_30_buffer [0:1];
  logic [63:0] PRED35_31_buffer [0:1];
  logic [63:0] PRED36_0_buffer [0:1];
  logic [63:0] PRED36_1_buffer [0:1];
  logic [63:0] PRED36_2_buffer [0:1];
  logic [63:0] PRED36_3_buffer [0:1];
  logic [63:0] PRED36_4_buffer [0:1];
  logic [63:0] PRED36_5_buffer [0:1];
  logic [63:0] PRED36_6_buffer [0:1];
  logic [63:0] PRED36_7_buffer [0:1];
  logic [63:0] PRED36_8_buffer [0:1];
  logic [63:0] PRED36_9_buffer [0:1];
  logic [63:0] PRED36_10_buffer [0:1];
  logic [63:0] PRED36_11_buffer [0:1];
  logic [63:0] PRED36_12_buffer [0:1];
  logic [63:0] PRED36_13_buffer [0:1];
  logic [63:0] PRED36_14_buffer [0:1];
  logic [63:0] PRED36_15_buffer [0:1];
  logic [63:0] PRED36_16_buffer [0:1];
  logic [63:0] PRED36_17_buffer [0:1];
  logic [63:0] PRED36_18_buffer [0:1];
  logic [63:0] PRED36_19_buffer [0:1];
  logic [63:0] PRED36_20_buffer [0:1];
  logic [63:0] PRED36_21_buffer [0:1];
  logic [63:0] PRED36_22_buffer [0:1];
  logic [63:0] PRED36_23_buffer [0:1];
  logic [63:0] PRED36_24_buffer [0:1];
  logic [63:0] PRED36_25_buffer [0:1];
  logic [63:0] PRED36_26_buffer [0:1];
  logic [63:0] PRED36_27_buffer [0:1];
  logic [63:0] PRED36_28_buffer [0:1];
  logic [63:0] PRED36_29_buffer [0:1];
  logic [63:0] PRED36_30_buffer [0:1];
  logic [63:0] PRED36_31_buffer [0:1];
  logic [63:0] PRED37_0_buffer [0:1];
  logic [63:0] PRED37_1_buffer [0:1];
  logic [63:0] PRED37_2_buffer [0:1];
  logic [63:0] PRED37_3_buffer [0:1];
  logic [63:0] PRED37_4_buffer [0:1];
  logic [63:0] PRED37_5_buffer [0:1];
  logic [63:0] PRED37_6_buffer [0:1];
  logic [63:0] PRED37_7_buffer [0:1];
  logic [63:0] PRED37_8_buffer [0:1];
  logic [63:0] PRED37_9_buffer [0:1];
  logic [63:0] PRED37_10_buffer [0:1];
  logic [63:0] PRED37_11_buffer [0:1];
  logic [63:0] PRED37_12_buffer [0:1];
  logic [63:0] PRED37_13_buffer [0:1];
  logic [63:0] PRED37_14_buffer [0:1];
  logic [63:0] PRED37_15_buffer [0:1];
  logic [63:0] PRED37_16_buffer [0:1];
  logic [63:0] PRED37_17_buffer [0:1];
  logic [63:0] PRED37_18_buffer [0:1];
  logic [63:0] PRED37_19_buffer [0:1];
  logic [63:0] PRED37_20_buffer [0:1];
  logic [63:0] PRED37_21_buffer [0:1];
  logic [63:0] PRED37_22_buffer [0:1];
  logic [63:0] PRED37_23_buffer [0:1];
  logic [63:0] PRED37_24_buffer [0:1];
  logic [63:0] PRED37_25_buffer [0:1];
  logic [63:0] PRED37_26_buffer [0:1];
  logic [63:0] PRED37_27_buffer [0:1];
  logic [63:0] PRED37_28_buffer [0:1];
  logic [63:0] PRED37_29_buffer [0:1];
  logic [63:0] PRED37_30_buffer [0:1];
  logic [63:0] PRED37_31_buffer [0:1];
  logic [63:0] PRED38_0_buffer [0:1];
  logic [63:0] PRED38_1_buffer [0:1];
  logic [63:0] PRED38_2_buffer [0:1];
  logic [63:0] PRED38_3_buffer [0:1];
  logic [63:0] PRED38_4_buffer [0:1];
  logic [63:0] PRED38_5_buffer [0:1];
  logic [63:0] PRED38_6_buffer [0:1];
  logic [63:0] PRED38_7_buffer [0:1];
  logic [63:0] PRED38_8_buffer [0:1];
  logic [63:0] PRED38_9_buffer [0:1];
  logic [63:0] PRED38_10_buffer [0:1];
  logic [63:0] PRED38_11_buffer [0:1];
  logic [63:0] PRED38_12_buffer [0:1];
  logic [63:0] PRED38_13_buffer [0:1];
  logic [63:0] PRED38_14_buffer [0:1];
  logic [63:0] PRED38_15_buffer [0:1];
  logic [63:0] PRED38_16_buffer [0:1];
  logic [63:0] PRED38_17_buffer [0:1];
  logic [63:0] PRED38_18_buffer [0:1];
  logic [63:0] PRED38_19_buffer [0:1];
  logic [63:0] PRED38_20_buffer [0:1];
  logic [63:0] PRED38_21_buffer [0:1];
  logic [63:0] PRED38_22_buffer [0:1];
  logic [63:0] PRED38_23_buffer [0:1];
  logic [63:0] PRED38_24_buffer [0:1];
  logic [63:0] PRED38_25_buffer [0:1];
  logic [63:0] PRED38_26_buffer [0:1];
  logic [63:0] PRED38_27_buffer [0:1];
  logic [63:0] PRED38_28_buffer [0:1];
  logic [63:0] PRED38_29_buffer [0:1];
  logic [63:0] PRED38_30_buffer [0:1];
  logic [63:0] PRED38_31_buffer [0:1];
  logic [63:0] PRED39_0_buffer [0:1];
  logic [63:0] PRED39_1_buffer [0:1];
  logic [63:0] PRED39_2_buffer [0:1];
  logic [63:0] PRED39_3_buffer [0:1];
  logic [63:0] PRED39_4_buffer [0:1];
  logic [63:0] PRED39_5_buffer [0:1];
  logic [63:0] PRED39_6_buffer [0:1];
  logic [63:0] PRED39_7_buffer [0:1];
  logic [63:0] PRED39_8_buffer [0:1];
  logic [63:0] PRED39_9_buffer [0:1];
  logic [63:0] PRED39_10_buffer [0:1];
  logic [63:0] PRED39_11_buffer [0:1];
  logic [63:0] PRED39_12_buffer [0:1];
  logic [63:0] PRED39_13_buffer [0:1];
  logic [63:0] PRED39_14_buffer [0:1];
  logic [63:0] PRED39_15_buffer [0:1];
  logic [63:0] PRED39_16_buffer [0:1];
  logic [63:0] PRED39_17_buffer [0:1];
  logic [63:0] PRED39_18_buffer [0:1];
  logic [63:0] PRED39_19_buffer [0:1];
  logic [63:0] PRED39_20_buffer [0:1];
  logic [63:0] PRED39_21_buffer [0:1];
  logic [63:0] PRED39_22_buffer [0:1];
  logic [63:0] PRED39_23_buffer [0:1];
  logic [63:0] PRED39_24_buffer [0:1];
  logic [63:0] PRED39_25_buffer [0:1];
  logic [63:0] PRED39_26_buffer [0:1];
  logic [63:0] PRED39_27_buffer [0:1];
  logic [63:0] PRED39_28_buffer [0:1];
  logic [63:0] PRED39_29_buffer [0:1];
  logic [63:0] PRED39_30_buffer [0:1];
  logic [63:0] PRED39_31_buffer [0:1];
  logic [63:0] PRED40_0_buffer [0:1];
  logic [63:0] PRED40_1_buffer [0:1];
  logic [63:0] PRED40_2_buffer [0:1];
  logic [63:0] PRED40_3_buffer [0:1];
  logic [63:0] PRED40_4_buffer [0:1];
  logic [63:0] PRED40_5_buffer [0:1];
  logic [63:0] PRED40_6_buffer [0:1];
  logic [63:0] PRED40_7_buffer [0:1];
  logic [63:0] PRED40_8_buffer [0:1];
  logic [63:0] PRED40_9_buffer [0:1];
  logic [63:0] PRED40_10_buffer [0:1];
  logic [63:0] PRED40_11_buffer [0:1];
  logic [63:0] PRED40_12_buffer [0:1];
  logic [63:0] PRED40_13_buffer [0:1];
  logic [63:0] PRED40_14_buffer [0:1];
  logic [63:0] PRED40_15_buffer [0:1];
  logic [63:0] PRED40_16_buffer [0:1];
  logic [63:0] PRED40_17_buffer [0:1];
  logic [63:0] PRED40_18_buffer [0:1];
  logic [63:0] PRED40_19_buffer [0:1];
  logic [63:0] PRED40_20_buffer [0:1];
  logic [63:0] PRED40_21_buffer [0:1];
  logic [63:0] PRED40_22_buffer [0:1];
  logic [63:0] PRED40_23_buffer [0:1];
  logic [63:0] PRED40_24_buffer [0:1];
  logic [63:0] PRED40_25_buffer [0:1];
  logic [63:0] PRED40_26_buffer [0:1];
  logic [63:0] PRED40_27_buffer [0:1];
  logic [63:0] PRED40_28_buffer [0:1];
  logic [63:0] PRED40_29_buffer [0:1];
  logic [63:0] PRED40_30_buffer [0:1];
  logic [63:0] PRED40_31_buffer [0:1];
  logic [63:0] PRED41_0_buffer [0:1];
  logic [63:0] PRED41_1_buffer [0:1];
  logic [63:0] PRED41_2_buffer [0:1];
  logic [63:0] PRED41_3_buffer [0:1];
  logic [63:0] PRED41_4_buffer [0:1];
  logic [63:0] PRED41_5_buffer [0:1];
  logic [63:0] PRED41_6_buffer [0:1];
  logic [63:0] PRED41_7_buffer [0:1];
  logic [63:0] PRED41_8_buffer [0:1];
  logic [63:0] PRED41_9_buffer [0:1];
  logic [63:0] PRED41_10_buffer [0:1];
  logic [63:0] PRED41_11_buffer [0:1];
  logic [63:0] PRED41_12_buffer [0:1];
  logic [63:0] PRED41_13_buffer [0:1];
  logic [63:0] PRED41_14_buffer [0:1];
  logic [63:0] PRED41_15_buffer [0:1];
  logic [63:0] PRED41_16_buffer [0:1];
  logic [63:0] PRED41_17_buffer [0:1];
  logic [63:0] PRED41_18_buffer [0:1];
  logic [63:0] PRED41_19_buffer [0:1];
  logic [63:0] PRED41_20_buffer [0:1];
  logic [63:0] PRED41_21_buffer [0:1];
  logic [63:0] PRED41_22_buffer [0:1];
  logic [63:0] PRED41_23_buffer [0:1];
  logic [63:0] PRED41_24_buffer [0:1];
  logic [63:0] PRED41_25_buffer [0:1];
  logic [63:0] PRED41_26_buffer [0:1];
  logic [63:0] PRED41_27_buffer [0:1];
  logic [63:0] PRED41_28_buffer [0:1];
  logic [63:0] PRED41_29_buffer [0:1];
  logic [63:0] PRED41_30_buffer [0:1];
  logic [63:0] PRED41_31_buffer [0:1];
  logic [63:0] PRED42_0_buffer [0:1];
  logic [63:0] PRED42_1_buffer [0:1];
  logic [63:0] PRED42_2_buffer [0:1];
  logic [63:0] PRED42_3_buffer [0:1];
  logic [63:0] PRED42_4_buffer [0:1];
  logic [63:0] PRED42_5_buffer [0:1];
  logic [63:0] PRED42_6_buffer [0:1];
  logic [63:0] PRED42_7_buffer [0:1];
  logic [63:0] PRED42_8_buffer [0:1];
  logic [63:0] PRED42_9_buffer [0:1];
  logic [63:0] PRED42_10_buffer [0:1];
  logic [63:0] PRED42_11_buffer [0:1];
  logic [63:0] PRED42_12_buffer [0:1];
  logic [63:0] PRED42_13_buffer [0:1];
  logic [63:0] PRED42_14_buffer [0:1];
  logic [63:0] PRED42_15_buffer [0:1];
  logic [63:0] PRED42_16_buffer [0:1];
  logic [63:0] PRED42_17_buffer [0:1];
  logic [63:0] PRED42_18_buffer [0:1];
  logic [63:0] PRED42_19_buffer [0:1];
  logic [63:0] PRED42_20_buffer [0:1];
  logic [63:0] PRED42_21_buffer [0:1];
  logic [63:0] PRED42_22_buffer [0:1];
  logic [63:0] PRED42_23_buffer [0:1];
  logic [63:0] PRED42_24_buffer [0:1];
  logic [63:0] PRED42_25_buffer [0:1];
  logic [63:0] PRED42_26_buffer [0:1];
  logic [63:0] PRED42_27_buffer [0:1];
  logic [63:0] PRED42_28_buffer [0:1];
  logic [63:0] PRED42_29_buffer [0:1];
  logic [63:0] PRED42_30_buffer [0:1];
  logic [63:0] PRED42_31_buffer [0:1];
  logic [63:0] PRED43_0_buffer [0:1];
  logic [63:0] PRED43_1_buffer [0:1];
  logic [63:0] PRED43_2_buffer [0:1];
  logic [63:0] PRED43_3_buffer [0:1];
  logic [63:0] PRED43_4_buffer [0:1];
  logic [63:0] PRED43_5_buffer [0:1];
  logic [63:0] PRED43_6_buffer [0:1];
  logic [63:0] PRED43_7_buffer [0:1];
  logic [63:0] PRED43_8_buffer [0:1];
  logic [63:0] PRED43_9_buffer [0:1];
  logic [63:0] PRED43_10_buffer [0:1];
  logic [63:0] PRED43_11_buffer [0:1];
  logic [63:0] PRED43_12_buffer [0:1];
  logic [63:0] PRED43_13_buffer [0:1];
  logic [63:0] PRED43_14_buffer [0:1];
  logic [63:0] PRED43_15_buffer [0:1];
  logic [63:0] PRED43_16_buffer [0:1];
  logic [63:0] PRED43_17_buffer [0:1];
  logic [63:0] PRED43_18_buffer [0:1];
  logic [63:0] PRED43_19_buffer [0:1];
  logic [63:0] PRED43_20_buffer [0:1];
  logic [63:0] PRED43_21_buffer [0:1];
  logic [63:0] PRED43_22_buffer [0:1];
  logic [63:0] PRED43_23_buffer [0:1];
  logic [63:0] PRED43_24_buffer [0:1];
  logic [63:0] PRED43_25_buffer [0:1];
  logic [63:0] PRED43_26_buffer [0:1];
  logic [63:0] PRED43_27_buffer [0:1];
  logic [63:0] PRED43_28_buffer [0:1];
  logic [63:0] PRED43_29_buffer [0:1];
  logic [63:0] PRED43_30_buffer [0:1];
  logic [63:0] PRED43_31_buffer [0:1];
  logic [63:0] PRED44_0_buffer [0:1];
  logic [63:0] PRED44_1_buffer [0:1];
  logic [63:0] PRED44_2_buffer [0:1];
  logic [63:0] PRED44_3_buffer [0:1];
  logic [63:0] PRED44_4_buffer [0:1];
  logic [63:0] PRED44_5_buffer [0:1];
  logic [63:0] PRED44_6_buffer [0:1];
  logic [63:0] PRED44_7_buffer [0:1];
  logic [63:0] PRED44_8_buffer [0:1];
  logic [63:0] PRED44_9_buffer [0:1];
  logic [63:0] PRED44_10_buffer [0:1];
  logic [63:0] PRED44_11_buffer [0:1];
  logic [63:0] PRED44_12_buffer [0:1];
  logic [63:0] PRED44_13_buffer [0:1];
  logic [63:0] PRED44_14_buffer [0:1];
  logic [63:0] PRED44_15_buffer [0:1];
  logic [63:0] PRED44_16_buffer [0:1];
  logic [63:0] PRED44_17_buffer [0:1];
  logic [63:0] PRED44_18_buffer [0:1];
  logic [63:0] PRED44_19_buffer [0:1];
  logic [63:0] PRED44_20_buffer [0:1];
  logic [63:0] PRED44_21_buffer [0:1];
  logic [63:0] PRED44_22_buffer [0:1];
  logic [63:0] PRED44_23_buffer [0:1];
  logic [63:0] PRED44_24_buffer [0:1];
  logic [63:0] PRED44_25_buffer [0:1];
  logic [63:0] PRED44_26_buffer [0:1];
  logic [63:0] PRED44_27_buffer [0:1];
  logic [63:0] PRED44_28_buffer [0:1];
  logic [63:0] PRED44_29_buffer [0:1];
  logic [63:0] PRED44_30_buffer [0:1];
  logic [63:0] PRED44_31_buffer [0:1];
  logic [63:0] PRED45_0_buffer [0:1];
  logic [63:0] PRED45_1_buffer [0:1];
  logic [63:0] PRED45_2_buffer [0:1];
  logic [63:0] PRED45_3_buffer [0:1];
  logic [63:0] PRED45_4_buffer [0:1];
  logic [63:0] PRED45_5_buffer [0:1];
  logic [63:0] PRED45_6_buffer [0:1];
  logic [63:0] PRED45_7_buffer [0:1];
  logic [63:0] PRED45_8_buffer [0:1];
  logic [63:0] PRED45_9_buffer [0:1];
  logic [63:0] PRED45_10_buffer [0:1];
  logic [63:0] PRED45_11_buffer [0:1];
  logic [63:0] PRED45_12_buffer [0:1];
  logic [63:0] PRED45_13_buffer [0:1];
  logic [63:0] PRED45_14_buffer [0:1];
  logic [63:0] PRED45_15_buffer [0:1];
  logic [63:0] PRED45_16_buffer [0:1];
  logic [63:0] PRED45_17_buffer [0:1];
  logic [63:0] PRED45_18_buffer [0:1];
  logic [63:0] PRED45_19_buffer [0:1];
  logic [63:0] PRED45_20_buffer [0:1];
  logic [63:0] PRED45_21_buffer [0:1];
  logic [63:0] PRED45_22_buffer [0:1];
  logic [63:0] PRED45_23_buffer [0:1];
  logic [63:0] PRED45_24_buffer [0:1];
  logic [63:0] PRED45_25_buffer [0:1];
  logic [63:0] PRED45_26_buffer [0:1];
  logic [63:0] PRED45_27_buffer [0:1];
  logic [63:0] PRED45_28_buffer [0:1];
  logic [63:0] PRED45_29_buffer [0:1];
  logic [63:0] PRED45_30_buffer [0:1];
  logic [63:0] PRED45_31_buffer [0:1];
  logic [63:0] PRED46_0_buffer [0:1];
  logic [63:0] PRED46_1_buffer [0:1];
  logic [63:0] PRED46_2_buffer [0:1];
  logic [63:0] PRED46_3_buffer [0:1];
  logic [63:0] PRED46_4_buffer [0:1];
  logic [63:0] PRED46_5_buffer [0:1];
  logic [63:0] PRED46_6_buffer [0:1];
  logic [63:0] PRED46_7_buffer [0:1];
  logic [63:0] PRED46_8_buffer [0:1];
  logic [63:0] PRED46_9_buffer [0:1];
  logic [63:0] PRED46_10_buffer [0:1];
  logic [63:0] PRED46_11_buffer [0:1];
  logic [63:0] PRED46_12_buffer [0:1];
  logic [63:0] PRED46_13_buffer [0:1];
  logic [63:0] PRED46_14_buffer [0:1];
  logic [63:0] PRED46_15_buffer [0:1];
  logic [63:0] PRED46_16_buffer [0:1];
  logic [63:0] PRED46_17_buffer [0:1];
  logic [63:0] PRED46_18_buffer [0:1];
  logic [63:0] PRED46_19_buffer [0:1];
  logic [63:0] PRED46_20_buffer [0:1];
  logic [63:0] PRED46_21_buffer [0:1];
  logic [63:0] PRED46_22_buffer [0:1];
  logic [63:0] PRED46_23_buffer [0:1];
  logic [63:0] PRED46_24_buffer [0:1];
  logic [63:0] PRED46_25_buffer [0:1];
  logic [63:0] PRED46_26_buffer [0:1];
  logic [63:0] PRED46_27_buffer [0:1];
  logic [63:0] PRED46_28_buffer [0:1];
  logic [63:0] PRED46_29_buffer [0:1];
  logic [63:0] PRED46_30_buffer [0:1];
  logic [63:0] PRED46_31_buffer [0:1];
  logic [63:0] PRED47_0_buffer [0:1];
  logic [63:0] PRED47_1_buffer [0:1];
  logic [63:0] PRED47_2_buffer [0:1];
  logic [63:0] PRED47_3_buffer [0:1];
  logic [63:0] PRED47_4_buffer [0:1];
  logic [63:0] PRED47_5_buffer [0:1];
  logic [63:0] PRED47_6_buffer [0:1];
  logic [63:0] PRED47_7_buffer [0:1];
  logic [63:0] PRED47_8_buffer [0:1];
  logic [63:0] PRED47_9_buffer [0:1];
  logic [63:0] PRED47_10_buffer [0:1];
  logic [63:0] PRED47_11_buffer [0:1];
  logic [63:0] PRED47_12_buffer [0:1];
  logic [63:0] PRED47_13_buffer [0:1];
  logic [63:0] PRED47_14_buffer [0:1];
  logic [63:0] PRED47_15_buffer [0:1];
  logic [63:0] PRED47_16_buffer [0:1];
  logic [63:0] PRED47_17_buffer [0:1];
  logic [63:0] PRED47_18_buffer [0:1];
  logic [63:0] PRED47_19_buffer [0:1];
  logic [63:0] PRED47_20_buffer [0:1];
  logic [63:0] PRED47_21_buffer [0:1];
  logic [63:0] PRED47_22_buffer [0:1];
  logic [63:0] PRED47_23_buffer [0:1];
  logic [63:0] PRED47_24_buffer [0:1];
  logic [63:0] PRED47_25_buffer [0:1];
  logic [63:0] PRED47_26_buffer [0:1];
  logic [63:0] PRED47_27_buffer [0:1];
  logic [63:0] PRED47_28_buffer [0:1];
  logic [63:0] PRED47_29_buffer [0:1];
  logic [63:0] PRED47_30_buffer [0:1];
  logic [63:0] PRED47_31_buffer [0:1];
  logic [63:0] PRED48_0_buffer [0:1];
  logic [63:0] PRED48_1_buffer [0:1];
  logic [63:0] PRED48_2_buffer [0:1];
  logic [63:0] PRED48_3_buffer [0:1];
  logic [63:0] PRED48_4_buffer [0:1];
  logic [63:0] PRED48_5_buffer [0:1];
  logic [63:0] PRED48_6_buffer [0:1];
  logic [63:0] PRED48_7_buffer [0:1];
  logic [63:0] PRED48_8_buffer [0:1];
  logic [63:0] PRED48_9_buffer [0:1];
  logic [63:0] PRED48_10_buffer [0:1];
  logic [63:0] PRED48_11_buffer [0:1];
  logic [63:0] PRED48_12_buffer [0:1];
  logic [63:0] PRED48_13_buffer [0:1];
  logic [63:0] PRED48_14_buffer [0:1];
  logic [63:0] PRED48_15_buffer [0:1];
  logic [63:0] PRED48_16_buffer [0:1];
  logic [63:0] PRED48_17_buffer [0:1];
  logic [63:0] PRED48_18_buffer [0:1];
  logic [63:0] PRED48_19_buffer [0:1];
  logic [63:0] PRED48_20_buffer [0:1];
  logic [63:0] PRED48_21_buffer [0:1];
  logic [63:0] PRED48_22_buffer [0:1];
  logic [63:0] PRED48_23_buffer [0:1];
  logic [63:0] PRED48_24_buffer [0:1];
  logic [63:0] PRED48_25_buffer [0:1];
  logic [63:0] PRED48_26_buffer [0:1];
  logic [63:0] PRED48_27_buffer [0:1];
  logic [63:0] PRED48_28_buffer [0:1];
  logic [63:0] PRED48_29_buffer [0:1];
  logic [63:0] PRED48_30_buffer [0:1];
  logic [63:0] PRED48_31_buffer [0:1];
  logic [63:0] PRED49_0_buffer [0:1];
  logic [63:0] PRED49_1_buffer [0:1];
  logic [63:0] PRED49_2_buffer [0:1];
  logic [63:0] PRED49_3_buffer [0:1];
  logic [63:0] PRED49_4_buffer [0:1];
  logic [63:0] PRED49_5_buffer [0:1];
  logic [63:0] PRED49_6_buffer [0:1];
  logic [63:0] PRED49_7_buffer [0:1];
  logic [63:0] PRED49_8_buffer [0:1];
  logic [63:0] PRED49_9_buffer [0:1];
  logic [63:0] PRED49_10_buffer [0:1];
  logic [63:0] PRED49_11_buffer [0:1];
  logic [63:0] PRED49_12_buffer [0:1];
  logic [63:0] PRED49_13_buffer [0:1];
  logic [63:0] PRED49_14_buffer [0:1];
  logic [63:0] PRED49_15_buffer [0:1];
  logic [63:0] PRED49_16_buffer [0:1];
  logic [63:0] PRED49_17_buffer [0:1];
  logic [63:0] PRED49_18_buffer [0:1];
  logic [63:0] PRED49_19_buffer [0:1];
  logic [63:0] PRED49_20_buffer [0:1];
  logic [63:0] PRED49_21_buffer [0:1];
  logic [63:0] PRED49_22_buffer [0:1];
  logic [63:0] PRED49_23_buffer [0:1];
  logic [63:0] PRED49_24_buffer [0:1];
  logic [63:0] PRED49_25_buffer [0:1];
  logic [63:0] PRED49_26_buffer [0:1];
  logic [63:0] PRED49_27_buffer [0:1];
  logic [63:0] PRED49_28_buffer [0:1];
  logic [63:0] PRED49_29_buffer [0:1];
  logic [63:0] PRED49_30_buffer [0:1];
  logic [63:0] PRED49_31_buffer [0:1];
  logic [63:0] PRED50_0_buffer [0:1];
  logic [63:0] PRED50_1_buffer [0:1];
  logic [63:0] PRED50_2_buffer [0:1];
  logic [63:0] PRED50_3_buffer [0:1];
  logic [63:0] PRED50_4_buffer [0:1];
  logic [63:0] PRED50_5_buffer [0:1];
  logic [63:0] PRED50_6_buffer [0:1];
  logic [63:0] PRED50_7_buffer [0:1];
  logic [63:0] PRED50_8_buffer [0:1];
  logic [63:0] PRED50_9_buffer [0:1];
  logic [63:0] PRED50_10_buffer [0:1];
  logic [63:0] PRED50_11_buffer [0:1];
  logic [63:0] PRED50_12_buffer [0:1];
  logic [63:0] PRED50_13_buffer [0:1];
  logic [63:0] PRED50_14_buffer [0:1];
  logic [63:0] PRED50_15_buffer [0:1];
  logic [63:0] PRED50_16_buffer [0:1];
  logic [63:0] PRED50_17_buffer [0:1];
  logic [63:0] PRED50_18_buffer [0:1];
  logic [63:0] PRED50_19_buffer [0:1];
  logic [63:0] PRED50_20_buffer [0:1];
  logic [63:0] PRED50_21_buffer [0:1];
  logic [63:0] PRED50_22_buffer [0:1];
  logic [63:0] PRED50_23_buffer [0:1];
  logic [63:0] PRED50_24_buffer [0:1];
  logic [63:0] PRED50_25_buffer [0:1];
  logic [63:0] PRED50_26_buffer [0:1];
  logic [63:0] PRED50_27_buffer [0:1];
  logic [63:0] PRED50_28_buffer [0:1];
  logic [63:0] PRED50_29_buffer [0:1];
  logic [63:0] PRED50_30_buffer [0:1];
  logic [63:0] PRED50_31_buffer [0:1];
  logic [63:0] PRED51_0_buffer [0:1];
  logic [63:0] PRED51_1_buffer [0:1];
  logic [63:0] PRED51_2_buffer [0:1];
  logic [63:0] PRED51_3_buffer [0:1];
  logic [63:0] PRED51_4_buffer [0:1];
  logic [63:0] PRED51_5_buffer [0:1];
  logic [63:0] PRED51_6_buffer [0:1];
  logic [63:0] PRED51_7_buffer [0:1];
  logic [63:0] PRED51_8_buffer [0:1];
  logic [63:0] PRED51_9_buffer [0:1];
  logic [63:0] PRED51_10_buffer [0:1];
  logic [63:0] PRED51_11_buffer [0:1];
  logic [63:0] PRED51_12_buffer [0:1];
  logic [63:0] PRED51_13_buffer [0:1];
  logic [63:0] PRED51_14_buffer [0:1];
  logic [63:0] PRED51_15_buffer [0:1];
  logic [63:0] PRED51_16_buffer [0:1];
  logic [63:0] PRED51_17_buffer [0:1];
  logic [63:0] PRED51_18_buffer [0:1];
  logic [63:0] PRED51_19_buffer [0:1];
  logic [63:0] PRED51_20_buffer [0:1];
  logic [63:0] PRED51_21_buffer [0:1];
  logic [63:0] PRED51_22_buffer [0:1];
  logic [63:0] PRED51_23_buffer [0:1];
  logic [63:0] PRED51_24_buffer [0:1];
  logic [63:0] PRED51_25_buffer [0:1];
  logic [63:0] PRED51_26_buffer [0:1];
  logic [63:0] PRED51_27_buffer [0:1];
  logic [63:0] PRED51_28_buffer [0:1];
  logic [63:0] PRED51_29_buffer [0:1];
  logic [63:0] PRED51_30_buffer [0:1];
  logic [63:0] PRED51_31_buffer [0:1];
  logic [63:0] PRED52_0_buffer [0:1];
  logic [63:0] PRED52_1_buffer [0:1];
  logic [63:0] PRED52_2_buffer [0:1];
  logic [63:0] PRED52_3_buffer [0:1];
  logic [63:0] PRED52_4_buffer [0:1];
  logic [63:0] PRED52_5_buffer [0:1];
  logic [63:0] PRED52_6_buffer [0:1];
  logic [63:0] PRED52_7_buffer [0:1];
  logic [63:0] PRED52_8_buffer [0:1];
  logic [63:0] PRED52_9_buffer [0:1];
  logic [63:0] PRED52_10_buffer [0:1];
  logic [63:0] PRED52_11_buffer [0:1];
  logic [63:0] PRED52_12_buffer [0:1];
  logic [63:0] PRED52_13_buffer [0:1];
  logic [63:0] PRED52_14_buffer [0:1];
  logic [63:0] PRED52_15_buffer [0:1];
  logic [63:0] PRED52_16_buffer [0:1];
  logic [63:0] PRED52_17_buffer [0:1];
  logic [63:0] PRED52_18_buffer [0:1];
  logic [63:0] PRED52_19_buffer [0:1];
  logic [63:0] PRED52_20_buffer [0:1];
  logic [63:0] PRED52_21_buffer [0:1];
  logic [63:0] PRED52_22_buffer [0:1];
  logic [63:0] PRED52_23_buffer [0:1];
  logic [63:0] PRED52_24_buffer [0:1];
  logic [63:0] PRED52_25_buffer [0:1];
  logic [63:0] PRED52_26_buffer [0:1];
  logic [63:0] PRED52_27_buffer [0:1];
  logic [63:0] PRED52_28_buffer [0:1];
  logic [63:0] PRED52_29_buffer [0:1];
  logic [63:0] PRED52_30_buffer [0:1];
  logic [63:0] PRED52_31_buffer [0:1];
  logic [63:0] PRED53_0_buffer [0:1];
  logic [63:0] PRED53_1_buffer [0:1];
  logic [63:0] PRED53_2_buffer [0:1];
  logic [63:0] PRED53_3_buffer [0:1];
  logic [63:0] PRED53_4_buffer [0:1];
  logic [63:0] PRED53_5_buffer [0:1];
  logic [63:0] PRED53_6_buffer [0:1];
  logic [63:0] PRED53_7_buffer [0:1];
  logic [63:0] PRED53_8_buffer [0:1];
  logic [63:0] PRED53_9_buffer [0:1];
  logic [63:0] PRED53_10_buffer [0:1];
  logic [63:0] PRED53_11_buffer [0:1];
  logic [63:0] PRED53_12_buffer [0:1];
  logic [63:0] PRED53_13_buffer [0:1];
  logic [63:0] PRED53_14_buffer [0:1];
  logic [63:0] PRED53_15_buffer [0:1];
  logic [63:0] PRED53_16_buffer [0:1];
  logic [63:0] PRED53_17_buffer [0:1];
  logic [63:0] PRED53_18_buffer [0:1];
  logic [63:0] PRED53_19_buffer [0:1];
  logic [63:0] PRED53_20_buffer [0:1];
  logic [63:0] PRED53_21_buffer [0:1];
  logic [63:0] PRED53_22_buffer [0:1];
  logic [63:0] PRED53_23_buffer [0:1];
  logic [63:0] PRED53_24_buffer [0:1];
  logic [63:0] PRED53_25_buffer [0:1];
  logic [63:0] PRED53_26_buffer [0:1];
  logic [63:0] PRED53_27_buffer [0:1];
  logic [63:0] PRED53_28_buffer [0:1];
  logic [63:0] PRED53_29_buffer [0:1];
  logic [63:0] PRED53_30_buffer [0:1];
  logic [63:0] PRED53_31_buffer [0:1];
  logic [63:0] PRED54_0_buffer [0:1];
  logic [63:0] PRED54_1_buffer [0:1];
  logic [63:0] PRED54_2_buffer [0:1];
  logic [63:0] PRED54_3_buffer [0:1];
  logic [63:0] PRED54_4_buffer [0:1];
  logic [63:0] PRED54_5_buffer [0:1];
  logic [63:0] PRED54_6_buffer [0:1];
  logic [63:0] PRED54_7_buffer [0:1];
  logic [63:0] PRED54_8_buffer [0:1];
  logic [63:0] PRED54_9_buffer [0:1];
  logic [63:0] PRED54_10_buffer [0:1];
  logic [63:0] PRED54_11_buffer [0:1];
  logic [63:0] PRED54_12_buffer [0:1];
  logic [63:0] PRED54_13_buffer [0:1];
  logic [63:0] PRED54_14_buffer [0:1];
  logic [63:0] PRED54_15_buffer [0:1];
  logic [63:0] PRED54_16_buffer [0:1];
  logic [63:0] PRED54_17_buffer [0:1];
  logic [63:0] PRED54_18_buffer [0:1];
  logic [63:0] PRED54_19_buffer [0:1];
  logic [63:0] PRED54_20_buffer [0:1];
  logic [63:0] PRED54_21_buffer [0:1];
  logic [63:0] PRED54_22_buffer [0:1];
  logic [63:0] PRED54_23_buffer [0:1];
  logic [63:0] PRED54_24_buffer [0:1];
  logic [63:0] PRED54_25_buffer [0:1];
  logic [63:0] PRED54_26_buffer [0:1];
  logic [63:0] PRED54_27_buffer [0:1];
  logic [63:0] PRED54_28_buffer [0:1];
  logic [63:0] PRED54_29_buffer [0:1];
  logic [63:0] PRED54_30_buffer [0:1];
  logic [63:0] PRED54_31_buffer [0:1];
  logic [63:0] PRED55_0_buffer [0:1];
  logic [63:0] PRED55_1_buffer [0:1];
  logic [63:0] PRED55_2_buffer [0:1];
  logic [63:0] PRED55_3_buffer [0:1];
  logic [63:0] PRED55_4_buffer [0:1];
  logic [63:0] PRED55_5_buffer [0:1];
  logic [63:0] PRED55_6_buffer [0:1];
  logic [63:0] PRED55_7_buffer [0:1];
  logic [63:0] PRED55_8_buffer [0:1];
  logic [63:0] PRED55_9_buffer [0:1];
  logic [63:0] PRED55_10_buffer [0:1];
  logic [63:0] PRED55_11_buffer [0:1];
  logic [63:0] PRED55_12_buffer [0:1];
  logic [63:0] PRED55_13_buffer [0:1];
  logic [63:0] PRED55_14_buffer [0:1];
  logic [63:0] PRED55_15_buffer [0:1];
  logic [63:0] PRED55_16_buffer [0:1];
  logic [63:0] PRED55_17_buffer [0:1];
  logic [63:0] PRED55_18_buffer [0:1];
  logic [63:0] PRED55_19_buffer [0:1];
  logic [63:0] PRED55_20_buffer [0:1];
  logic [63:0] PRED55_21_buffer [0:1];
  logic [63:0] PRED55_22_buffer [0:1];
  logic [63:0] PRED55_23_buffer [0:1];
  logic [63:0] PRED55_24_buffer [0:1];
  logic [63:0] PRED55_25_buffer [0:1];
  logic [63:0] PRED55_26_buffer [0:1];
  logic [63:0] PRED55_27_buffer [0:1];
  logic [63:0] PRED55_28_buffer [0:1];
  logic [63:0] PRED55_29_buffer [0:1];
  logic [63:0] PRED55_30_buffer [0:1];
  logic [63:0] PRED55_31_buffer [0:1];
  logic [63:0] PRED56_0_buffer [0:1];
  logic [63:0] PRED56_1_buffer [0:1];
  logic [63:0] PRED56_2_buffer [0:1];
  logic [63:0] PRED56_3_buffer [0:1];
  logic [63:0] PRED56_4_buffer [0:1];
  logic [63:0] PRED56_5_buffer [0:1];
  logic [63:0] PRED56_6_buffer [0:1];
  logic [63:0] PRED56_7_buffer [0:1];
  logic [63:0] PRED56_8_buffer [0:1];
  logic [63:0] PRED56_9_buffer [0:1];
  logic [63:0] PRED56_10_buffer [0:1];
  logic [63:0] PRED56_11_buffer [0:1];
  logic [63:0] PRED56_12_buffer [0:1];
  logic [63:0] PRED56_13_buffer [0:1];
  logic [63:0] PRED56_14_buffer [0:1];
  logic [63:0] PRED56_15_buffer [0:1];
  logic [63:0] PRED56_16_buffer [0:1];
  logic [63:0] PRED56_17_buffer [0:1];
  logic [63:0] PRED56_18_buffer [0:1];
  logic [63:0] PRED56_19_buffer [0:1];
  logic [63:0] PRED56_20_buffer [0:1];
  logic [63:0] PRED56_21_buffer [0:1];
  logic [63:0] PRED56_22_buffer [0:1];
  logic [63:0] PRED56_23_buffer [0:1];
  logic [63:0] PRED56_24_buffer [0:1];
  logic [63:0] PRED56_25_buffer [0:1];
  logic [63:0] PRED56_26_buffer [0:1];
  logic [63:0] PRED56_27_buffer [0:1];
  logic [63:0] PRED56_28_buffer [0:1];
  logic [63:0] PRED56_29_buffer [0:1];
  logic [63:0] PRED56_30_buffer [0:1];
  logic [63:0] PRED56_31_buffer [0:1];
  logic [63:0] PRED57_0_buffer [0:1];
  logic [63:0] PRED57_1_buffer [0:1];
  logic [63:0] PRED57_2_buffer [0:1];
  logic [63:0] PRED57_3_buffer [0:1];
  logic [63:0] PRED57_4_buffer [0:1];
  logic [63:0] PRED57_5_buffer [0:1];
  logic [63:0] PRED57_6_buffer [0:1];
  logic [63:0] PRED57_7_buffer [0:1];
  logic [63:0] PRED57_8_buffer [0:1];
  logic [63:0] PRED57_9_buffer [0:1];
  logic [63:0] PRED57_10_buffer [0:1];
  logic [63:0] PRED57_11_buffer [0:1];
  logic [63:0] PRED57_12_buffer [0:1];
  logic [63:0] PRED57_13_buffer [0:1];
  logic [63:0] PRED57_14_buffer [0:1];
  logic [63:0] PRED57_15_buffer [0:1];
  logic [63:0] PRED57_16_buffer [0:1];
  logic [63:0] PRED57_17_buffer [0:1];
  logic [63:0] PRED57_18_buffer [0:1];
  logic [63:0] PRED57_19_buffer [0:1];
  logic [63:0] PRED57_20_buffer [0:1];
  logic [63:0] PRED57_21_buffer [0:1];
  logic [63:0] PRED57_22_buffer [0:1];
  logic [63:0] PRED57_23_buffer [0:1];
  logic [63:0] PRED57_24_buffer [0:1];
  logic [63:0] PRED57_25_buffer [0:1];
  logic [63:0] PRED57_26_buffer [0:1];
  logic [63:0] PRED57_27_buffer [0:1];
  logic [63:0] PRED57_28_buffer [0:1];
  logic [63:0] PRED57_29_buffer [0:1];
  logic [63:0] PRED57_30_buffer [0:1];
  logic [63:0] PRED57_31_buffer [0:1];
  logic [63:0] PRED58_0_buffer [0:1];
  logic [63:0] PRED58_1_buffer [0:1];
  logic [63:0] PRED58_2_buffer [0:1];
  logic [63:0] PRED58_3_buffer [0:1];
  logic [63:0] PRED58_4_buffer [0:1];
  logic [63:0] PRED58_5_buffer [0:1];
  logic [63:0] PRED58_6_buffer [0:1];
  logic [63:0] PRED58_7_buffer [0:1];
  logic [63:0] PRED58_8_buffer [0:1];
  logic [63:0] PRED58_9_buffer [0:1];
  logic [63:0] PRED58_10_buffer [0:1];
  logic [63:0] PRED58_11_buffer [0:1];
  logic [63:0] PRED58_12_buffer [0:1];
  logic [63:0] PRED58_13_buffer [0:1];
  logic [63:0] PRED58_14_buffer [0:1];
  logic [63:0] PRED58_15_buffer [0:1];
  logic [63:0] PRED58_16_buffer [0:1];
  logic [63:0] PRED58_17_buffer [0:1];
  logic [63:0] PRED58_18_buffer [0:1];
  logic [63:0] PRED58_19_buffer [0:1];
  logic [63:0] PRED58_20_buffer [0:1];
  logic [63:0] PRED58_21_buffer [0:1];
  logic [63:0] PRED58_22_buffer [0:1];
  logic [63:0] PRED58_23_buffer [0:1];
  logic [63:0] PRED58_24_buffer [0:1];
  logic [63:0] PRED58_25_buffer [0:1];
  logic [63:0] PRED58_26_buffer [0:1];
  logic [63:0] PRED58_27_buffer [0:1];
  logic [63:0] PRED58_28_buffer [0:1];
  logic [63:0] PRED58_29_buffer [0:1];
  logic [63:0] PRED58_30_buffer [0:1];
  logic [63:0] PRED58_31_buffer [0:1];
  logic [63:0] PRED59_0_buffer [0:1];
  logic [63:0] PRED59_1_buffer [0:1];
  logic [63:0] PRED59_2_buffer [0:1];
  logic [63:0] PRED59_3_buffer [0:1];
  logic [63:0] PRED59_4_buffer [0:1];
  logic [63:0] PRED59_5_buffer [0:1];
  logic [63:0] PRED59_6_buffer [0:1];
  logic [63:0] PRED59_7_buffer [0:1];
  logic [63:0] PRED59_8_buffer [0:1];
  logic [63:0] PRED59_9_buffer [0:1];
  logic [63:0] PRED59_10_buffer [0:1];
  logic [63:0] PRED59_11_buffer [0:1];
  logic [63:0] PRED59_12_buffer [0:1];
  logic [63:0] PRED59_13_buffer [0:1];
  logic [63:0] PRED59_14_buffer [0:1];
  logic [63:0] PRED59_15_buffer [0:1];
  logic [63:0] PRED59_16_buffer [0:1];
  logic [63:0] PRED59_17_buffer [0:1];
  logic [63:0] PRED59_18_buffer [0:1];
  logic [63:0] PRED59_19_buffer [0:1];
  logic [63:0] PRED59_20_buffer [0:1];
  logic [63:0] PRED59_21_buffer [0:1];
  logic [63:0] PRED59_22_buffer [0:1];
  logic [63:0] PRED59_23_buffer [0:1];
  logic [63:0] PRED59_24_buffer [0:1];
  logic [63:0] PRED59_25_buffer [0:1];
  logic [63:0] PRED59_26_buffer [0:1];
  logic [63:0] PRED59_27_buffer [0:1];
  logic [63:0] PRED59_28_buffer [0:1];
  logic [63:0] PRED59_29_buffer [0:1];
  logic [63:0] PRED59_30_buffer [0:1];
  logic [63:0] PRED59_31_buffer [0:1];
  logic [63:0] PRED60_0_buffer [0:1];
  logic [63:0] PRED60_1_buffer [0:1];
  logic [63:0] PRED60_2_buffer [0:1];
  logic [63:0] PRED60_3_buffer [0:1];
  logic [63:0] PRED60_4_buffer [0:1];
  logic [63:0] PRED60_5_buffer [0:1];
  logic [63:0] PRED60_6_buffer [0:1];
  logic [63:0] PRED60_7_buffer [0:1];
  logic [63:0] PRED60_8_buffer [0:1];
  logic [63:0] PRED60_9_buffer [0:1];
  logic [63:0] PRED60_10_buffer [0:1];
  logic [63:0] PRED60_11_buffer [0:1];
  logic [63:0] PRED60_12_buffer [0:1];
  logic [63:0] PRED60_13_buffer [0:1];
  logic [63:0] PRED60_14_buffer [0:1];
  logic [63:0] PRED60_15_buffer [0:1];
  logic [63:0] PRED60_16_buffer [0:1];
  logic [63:0] PRED60_17_buffer [0:1];
  logic [63:0] PRED60_18_buffer [0:1];
  logic [63:0] PRED60_19_buffer [0:1];
  logic [63:0] PRED60_20_buffer [0:1];
  logic [63:0] PRED60_21_buffer [0:1];
  logic [63:0] PRED60_22_buffer [0:1];
  logic [63:0] PRED60_23_buffer [0:1];
  logic [63:0] PRED60_24_buffer [0:1];
  logic [63:0] PRED60_25_buffer [0:1];
  logic [63:0] PRED60_26_buffer [0:1];
  logic [63:0] PRED60_27_buffer [0:1];
  logic [63:0] PRED60_28_buffer [0:1];
  logic [63:0] PRED60_29_buffer [0:1];
  logic [63:0] PRED60_30_buffer [0:1];
  logic [63:0] PRED60_31_buffer [0:1];
  logic [63:0] PRED61_0_buffer [0:1];
  logic [63:0] PRED61_1_buffer [0:1];
  logic [63:0] PRED61_2_buffer [0:1];
  logic [63:0] PRED61_3_buffer [0:1];
  logic [63:0] PRED61_4_buffer [0:1];
  logic [63:0] PRED61_5_buffer [0:1];
  logic [63:0] PRED61_6_buffer [0:1];
  logic [63:0] PRED61_7_buffer [0:1];
  logic [63:0] PRED61_8_buffer [0:1];
  logic [63:0] PRED61_9_buffer [0:1];
  logic [63:0] PRED61_10_buffer [0:1];
  logic [63:0] PRED61_11_buffer [0:1];
  logic [63:0] PRED61_12_buffer [0:1];
  logic [63:0] PRED61_13_buffer [0:1];
  logic [63:0] PRED61_14_buffer [0:1];
  logic [63:0] PRED61_15_buffer [0:1];
  logic [63:0] PRED61_16_buffer [0:1];
  logic [63:0] PRED61_17_buffer [0:1];
  logic [63:0] PRED61_18_buffer [0:1];
  logic [63:0] PRED61_19_buffer [0:1];
  logic [63:0] PRED61_20_buffer [0:1];
  logic [63:0] PRED61_21_buffer [0:1];
  logic [63:0] PRED61_22_buffer [0:1];
  logic [63:0] PRED61_23_buffer [0:1];
  logic [63:0] PRED61_24_buffer [0:1];
  logic [63:0] PRED61_25_buffer [0:1];
  logic [63:0] PRED61_26_buffer [0:1];
  logic [63:0] PRED61_27_buffer [0:1];
  logic [63:0] PRED61_28_buffer [0:1];
  logic [63:0] PRED61_29_buffer [0:1];
  logic [63:0] PRED61_30_buffer [0:1];
  logic [63:0] PRED61_31_buffer [0:1];
  logic [63:0] PRED62_0_buffer [0:1];
  logic [63:0] PRED62_1_buffer [0:1];
  logic [63:0] PRED62_2_buffer [0:1];
  logic [63:0] PRED62_3_buffer [0:1];
  logic [63:0] PRED62_4_buffer [0:1];
  logic [63:0] PRED62_5_buffer [0:1];
  logic [63:0] PRED62_6_buffer [0:1];
  logic [63:0] PRED62_7_buffer [0:1];
  logic [63:0] PRED62_8_buffer [0:1];
  logic [63:0] PRED62_9_buffer [0:1];
  logic [63:0] PRED62_10_buffer [0:1];
  logic [63:0] PRED62_11_buffer [0:1];
  logic [63:0] PRED62_12_buffer [0:1];
  logic [63:0] PRED62_13_buffer [0:1];
  logic [63:0] PRED62_14_buffer [0:1];
  logic [63:0] PRED62_15_buffer [0:1];
  logic [63:0] PRED62_16_buffer [0:1];
  logic [63:0] PRED62_17_buffer [0:1];
  logic [63:0] PRED62_18_buffer [0:1];
  logic [63:0] PRED62_19_buffer [0:1];
  logic [63:0] PRED62_20_buffer [0:1];
  logic [63:0] PRED62_21_buffer [0:1];
  logic [63:0] PRED62_22_buffer [0:1];
  logic [63:0] PRED62_23_buffer [0:1];
  logic [63:0] PRED62_24_buffer [0:1];
  logic [63:0] PRED62_25_buffer [0:1];
  logic [63:0] PRED62_26_buffer [0:1];
  logic [63:0] PRED62_27_buffer [0:1];
  logic [63:0] PRED62_28_buffer [0:1];
  logic [63:0] PRED62_29_buffer [0:1];
  logic [63:0] PRED62_30_buffer [0:1];
  logic [63:0] PRED62_31_buffer [0:1];
  logic [63:0] PRED63_0_buffer [0:1];
  logic [63:0] PRED63_1_buffer [0:1];
  logic [63:0] PRED63_2_buffer [0:1];
  logic [63:0] PRED63_3_buffer [0:1];
  logic [63:0] PRED63_4_buffer [0:1];
  logic [63:0] PRED63_5_buffer [0:1];
  logic [63:0] PRED63_6_buffer [0:1];
  logic [63:0] PRED63_7_buffer [0:1];
  logic [63:0] PRED63_8_buffer [0:1];
  logic [63:0] PRED63_9_buffer [0:1];
  logic [63:0] PRED63_10_buffer [0:1];
  logic [63:0] PRED63_11_buffer [0:1];
  logic [63:0] PRED63_12_buffer [0:1];
  logic [63:0] PRED63_13_buffer [0:1];
  logic [63:0] PRED63_14_buffer [0:1];
  logic [63:0] PRED63_15_buffer [0:1];
  logic [63:0] PRED63_16_buffer [0:1];
  logic [63:0] PRED63_17_buffer [0:1];
  logic [63:0] PRED63_18_buffer [0:1];
  logic [63:0] PRED63_19_buffer [0:1];
  logic [63:0] PRED63_20_buffer [0:1];
  logic [63:0] PRED63_21_buffer [0:1];
  logic [63:0] PRED63_22_buffer [0:1];
  logic [63:0] PRED63_23_buffer [0:1];
  logic [63:0] PRED63_24_buffer [0:1];
  logic [63:0] PRED63_25_buffer [0:1];
  logic [63:0] PRED63_26_buffer [0:1];
  logic [63:0] PRED63_27_buffer [0:1];
  logic [63:0] PRED63_28_buffer [0:1];
  logic [63:0] PRED63_29_buffer [0:1];
  logic [63:0] PRED63_30_buffer [0:1];
  logic [63:0] PRED63_31_buffer [0:1];

  // initiate warp signals (1 if there is a change in one of the buffers)
  logic warp0_sig;
  logic warp1_sig;
  logic warp2_sig;
  logic warp3_sig;
  logic warp4_sig;
  logic warp5_sig;
  logic warp6_sig;
  logic warp7_sig;


  // Initialize the output tracker file
  initial begin
    f = $fopen("h_tracker_pred.txt", "w");
    $fwrite(f, "=====================================================\n");
    $fwrite(f, "              Harmonica Tracker v1");
    $fwrite(f, " \n=====================================================\n\n");

  end


  // Need to differentiate between different warps time instruction and changes to memory and registers

  // Put information into the buffer // FIXME, code bloat // for loop  -- syntax for printing is not correct, so i just copied and paste from C++ code // FIXME
  always @ (edge clk) begin
    PRED0_0_buffer[clk] = PRED0[0];
    PRED0_1_buffer[clk] = PRED0[1];
    PRED0_2_buffer[clk] = PRED0[2];
    PRED0_3_buffer[clk] = PRED0[3];
    PRED0_4_buffer[clk] = PRED0[4];
    PRED0_5_buffer[clk] = PRED0[5];
    PRED0_6_buffer[clk] = PRED0[6];
    PRED0_7_buffer[clk] = PRED0[7];
    PRED0_8_buffer[clk] = PRED0[8];
    PRED0_9_buffer[clk] = PRED0[9];
    PRED0_10_buffer[clk] = PRED0[10];
    PRED0_11_buffer[clk] = PRED0[11];
    PRED0_12_buffer[clk] = PRED0[12];
    PRED0_13_buffer[clk] = PRED0[13];
    PRED0_14_buffer[clk] = PRED0[14];
    PRED0_15_buffer[clk] = PRED0[15];
    PRED0_16_buffer[clk] = PRED0[16];
    PRED0_17_buffer[clk] = PRED0[17];
    PRED0_18_buffer[clk] = PRED0[18];
    PRED0_19_buffer[clk] = PRED0[19];
    PRED0_20_buffer[clk] = PRED0[20];
    PRED0_21_buffer[clk] = PRED0[21];
    PRED0_22_buffer[clk] = PRED0[22];
    PRED0_23_buffer[clk] = PRED0[23];
    PRED0_24_buffer[clk] = PRED0[24];
    PRED0_25_buffer[clk] = PRED0[25];
    PRED0_26_buffer[clk] = PRED0[26];
    PRED0_27_buffer[clk] = PRED0[27];
    PRED0_28_buffer[clk] = PRED0[28];
    PRED0_29_buffer[clk] = PRED0[29];
    PRED0_30_buffer[clk] = PRED0[30];
    PRED0_31_buffer[clk] = PRED0[31];
    PRED1_0_buffer[clk] = PRED1[0];
    PRED1_1_buffer[clk] = PRED1[1];
    PRED1_2_buffer[clk] = PRED1[2];
    PRED1_3_buffer[clk] = PRED1[3];
    PRED1_4_buffer[clk] = PRED1[4];
    PRED1_5_buffer[clk] = PRED1[5];
    PRED1_6_buffer[clk] = PRED1[6];
    PRED1_7_buffer[clk] = PRED1[7];
    PRED1_8_buffer[clk] = PRED1[8];
    PRED1_9_buffer[clk] = PRED1[9];
    PRED1_10_buffer[clk] = PRED1[10];
    PRED1_11_buffer[clk] = PRED1[11];
    PRED1_12_buffer[clk] = PRED1[12];
    PRED1_13_buffer[clk] = PRED1[13];
    PRED1_14_buffer[clk] = PRED1[14];
    PRED1_15_buffer[clk] = PRED1[15];
    PRED1_16_buffer[clk] = PRED1[16];
    PRED1_17_buffer[clk] = PRED1[17];
    PRED1_18_buffer[clk] = PRED1[18];
    PRED1_19_buffer[clk] = PRED1[19];
    PRED1_20_buffer[clk] = PRED1[20];
    PRED1_21_buffer[clk] = PRED1[21];
    PRED1_22_buffer[clk] = PRED1[22];
    PRED1_23_buffer[clk] = PRED1[23];
    PRED1_24_buffer[clk] = PRED1[24];
    PRED1_25_buffer[clk] = PRED1[25];
    PRED1_26_buffer[clk] = PRED1[26];
    PRED1_27_buffer[clk] = PRED1[27];
    PRED1_28_buffer[clk] = PRED1[28];
    PRED1_29_buffer[clk] = PRED1[29];
    PRED1_30_buffer[clk] = PRED1[30];
    PRED1_31_buffer[clk] = PRED1[31];
    PRED2_0_buffer[clk] = PRED2[0];
    PRED2_1_buffer[clk] = PRED2[1];
    PRED2_2_buffer[clk] = PRED2[2];
    PRED2_3_buffer[clk] = PRED2[3];
    PRED2_4_buffer[clk] = PRED2[4];
    PRED2_5_buffer[clk] = PRED2[5];
    PRED2_6_buffer[clk] = PRED2[6];
    PRED2_7_buffer[clk] = PRED2[7];
    PRED2_8_buffer[clk] = PRED2[8];
    PRED2_9_buffer[clk] = PRED2[9];
    PRED2_10_buffer[clk] = PRED2[10];
    PRED2_11_buffer[clk] = PRED2[11];
    PRED2_12_buffer[clk] = PRED2[12];
    PRED2_13_buffer[clk] = PRED2[13];
    PRED2_14_buffer[clk] = PRED2[14];
    PRED2_15_buffer[clk] = PRED2[15];
    PRED2_16_buffer[clk] = PRED2[16];
    PRED2_17_buffer[clk] = PRED2[17];
    PRED2_18_buffer[clk] = PRED2[18];
    PRED2_19_buffer[clk] = PRED2[19];
    PRED2_20_buffer[clk] = PRED2[20];
    PRED2_21_buffer[clk] = PRED2[21];
    PRED2_22_buffer[clk] = PRED2[22];
    PRED2_23_buffer[clk] = PRED2[23];
    PRED2_24_buffer[clk] = PRED2[24];
    PRED2_25_buffer[clk] = PRED2[25];
    PRED2_26_buffer[clk] = PRED2[26];
    PRED2_27_buffer[clk] = PRED2[27];
    PRED2_28_buffer[clk] = PRED2[28];
    PRED2_29_buffer[clk] = PRED2[29];
    PRED2_30_buffer[clk] = PRED2[30];
    PRED2_31_buffer[clk] = PRED2[31];
    PRED3_0_buffer[clk] = PRED3[0];
    PRED3_1_buffer[clk] = PRED3[1];
    PRED3_2_buffer[clk] = PRED3[2];
    PRED3_3_buffer[clk] = PRED3[3];
    PRED3_4_buffer[clk] = PRED3[4];
    PRED3_5_buffer[clk] = PRED3[5];
    PRED3_6_buffer[clk] = PRED3[6];
    PRED3_7_buffer[clk] = PRED3[7];
    PRED3_8_buffer[clk] = PRED3[8];
    PRED3_9_buffer[clk] = PRED3[9];
    PRED3_10_buffer[clk] = PRED3[10];
    PRED3_11_buffer[clk] = PRED3[11];
    PRED3_12_buffer[clk] = PRED3[12];
    PRED3_13_buffer[clk] = PRED3[13];
    PRED3_14_buffer[clk] = PRED3[14];
    PRED3_15_buffer[clk] = PRED3[15];
    PRED3_16_buffer[clk] = PRED3[16];
    PRED3_17_buffer[clk] = PRED3[17];
    PRED3_18_buffer[clk] = PRED3[18];
    PRED3_19_buffer[clk] = PRED3[19];
    PRED3_20_buffer[clk] = PRED3[20];
    PRED3_21_buffer[clk] = PRED3[21];
    PRED3_22_buffer[clk] = PRED3[22];
    PRED3_23_buffer[clk] = PRED3[23];
    PRED3_24_buffer[clk] = PRED3[24];
    PRED3_25_buffer[clk] = PRED3[25];
    PRED3_26_buffer[clk] = PRED3[26];
    PRED3_27_buffer[clk] = PRED3[27];
    PRED3_28_buffer[clk] = PRED3[28];
    PRED3_29_buffer[clk] = PRED3[29];
    PRED3_30_buffer[clk] = PRED3[30];
    PRED3_31_buffer[clk] = PRED3[31];
    PRED4_0_buffer[clk] = PRED4[0];
    PRED4_1_buffer[clk] = PRED4[1];
    PRED4_2_buffer[clk] = PRED4[2];
    PRED4_3_buffer[clk] = PRED4[3];
    PRED4_4_buffer[clk] = PRED4[4];
    PRED4_5_buffer[clk] = PRED4[5];
    PRED4_6_buffer[clk] = PRED4[6];
    PRED4_7_buffer[clk] = PRED4[7];
    PRED4_8_buffer[clk] = PRED4[8];
    PRED4_9_buffer[clk] = PRED4[9];
    PRED4_10_buffer[clk] = PRED4[10];
    PRED4_11_buffer[clk] = PRED4[11];
    PRED4_12_buffer[clk] = PRED4[12];
    PRED4_13_buffer[clk] = PRED4[13];
    PRED4_14_buffer[clk] = PRED4[14];
    PRED4_15_buffer[clk] = PRED4[15];
    PRED4_16_buffer[clk] = PRED4[16];
    PRED4_17_buffer[clk] = PRED4[17];
    PRED4_18_buffer[clk] = PRED4[18];
    PRED4_19_buffer[clk] = PRED4[19];
    PRED4_20_buffer[clk] = PRED4[20];
    PRED4_21_buffer[clk] = PRED4[21];
    PRED4_22_buffer[clk] = PRED4[22];
    PRED4_23_buffer[clk] = PRED4[23];
    PRED4_24_buffer[clk] = PRED4[24];
    PRED4_25_buffer[clk] = PRED4[25];
    PRED4_26_buffer[clk] = PRED4[26];
    PRED4_27_buffer[clk] = PRED4[27];
    PRED4_28_buffer[clk] = PRED4[28];
    PRED4_29_buffer[clk] = PRED4[29];
    PRED4_30_buffer[clk] = PRED4[30];
    PRED4_31_buffer[clk] = PRED4[31];
    PRED5_0_buffer[clk] = PRED5[0];
    PRED5_1_buffer[clk] = PRED5[1];
    PRED5_2_buffer[clk] = PRED5[2];
    PRED5_3_buffer[clk] = PRED5[3];
    PRED5_4_buffer[clk] = PRED5[4];
    PRED5_5_buffer[clk] = PRED5[5];
    PRED5_6_buffer[clk] = PRED5[6];
    PRED5_7_buffer[clk] = PRED5[7];
    PRED5_8_buffer[clk] = PRED5[8];
    PRED5_9_buffer[clk] = PRED5[9];
    PRED5_10_buffer[clk] = PRED5[10];
    PRED5_11_buffer[clk] = PRED5[11];
    PRED5_12_buffer[clk] = PRED5[12];
    PRED5_13_buffer[clk] = PRED5[13];
    PRED5_14_buffer[clk] = PRED5[14];
    PRED5_15_buffer[clk] = PRED5[15];
    PRED5_16_buffer[clk] = PRED5[16];
    PRED5_17_buffer[clk] = PRED5[17];
    PRED5_18_buffer[clk] = PRED5[18];
    PRED5_19_buffer[clk] = PRED5[19];
    PRED5_20_buffer[clk] = PRED5[20];
    PRED5_21_buffer[clk] = PRED5[21];
    PRED5_22_buffer[clk] = PRED5[22];
    PRED5_23_buffer[clk] = PRED5[23];
    PRED5_24_buffer[clk] = PRED5[24];
    PRED5_25_buffer[clk] = PRED5[25];
    PRED5_26_buffer[clk] = PRED5[26];
    PRED5_27_buffer[clk] = PRED5[27];
    PRED5_28_buffer[clk] = PRED5[28];
    PRED5_29_buffer[clk] = PRED5[29];
    PRED5_30_buffer[clk] = PRED5[30];
    PRED5_31_buffer[clk] = PRED5[31];
    PRED6_0_buffer[clk] = PRED6[0];
    PRED6_1_buffer[clk] = PRED6[1];
    PRED6_2_buffer[clk] = PRED6[2];
    PRED6_3_buffer[clk] = PRED6[3];
    PRED6_4_buffer[clk] = PRED6[4];
    PRED6_5_buffer[clk] = PRED6[5];
    PRED6_6_buffer[clk] = PRED6[6];
    PRED6_7_buffer[clk] = PRED6[7];
    PRED6_8_buffer[clk] = PRED6[8];
    PRED6_9_buffer[clk] = PRED6[9];
    PRED6_10_buffer[clk] = PRED6[10];
    PRED6_11_buffer[clk] = PRED6[11];
    PRED6_12_buffer[clk] = PRED6[12];
    PRED6_13_buffer[clk] = PRED6[13];
    PRED6_14_buffer[clk] = PRED6[14];
    PRED6_15_buffer[clk] = PRED6[15];
    PRED6_16_buffer[clk] = PRED6[16];
    PRED6_17_buffer[clk] = PRED6[17];
    PRED6_18_buffer[clk] = PRED6[18];
    PRED6_19_buffer[clk] = PRED6[19];
    PRED6_20_buffer[clk] = PRED6[20];
    PRED6_21_buffer[clk] = PRED6[21];
    PRED6_22_buffer[clk] = PRED6[22];
    PRED6_23_buffer[clk] = PRED6[23];
    PRED6_24_buffer[clk] = PRED6[24];
    PRED6_25_buffer[clk] = PRED6[25];
    PRED6_26_buffer[clk] = PRED6[26];
    PRED6_27_buffer[clk] = PRED6[27];
    PRED6_28_buffer[clk] = PRED6[28];
    PRED6_29_buffer[clk] = PRED6[29];
    PRED6_30_buffer[clk] = PRED6[30];
    PRED6_31_buffer[clk] = PRED6[31];
    PRED7_0_buffer[clk] = PRED7[0];
    PRED7_1_buffer[clk] = PRED7[1];
    PRED7_2_buffer[clk] = PRED7[2];
    PRED7_3_buffer[clk] = PRED7[3];
    PRED7_4_buffer[clk] = PRED7[4];
    PRED7_5_buffer[clk] = PRED7[5];
    PRED7_6_buffer[clk] = PRED7[6];
    PRED7_7_buffer[clk] = PRED7[7];
    PRED7_8_buffer[clk] = PRED7[8];
    PRED7_9_buffer[clk] = PRED7[9];
    PRED7_10_buffer[clk] = PRED7[10];
    PRED7_11_buffer[clk] = PRED7[11];
    PRED7_12_buffer[clk] = PRED7[12];
    PRED7_13_buffer[clk] = PRED7[13];
    PRED7_14_buffer[clk] = PRED7[14];
    PRED7_15_buffer[clk] = PRED7[15];
    PRED7_16_buffer[clk] = PRED7[16];
    PRED7_17_buffer[clk] = PRED7[17];
    PRED7_18_buffer[clk] = PRED7[18];
    PRED7_19_buffer[clk] = PRED7[19];
    PRED7_20_buffer[clk] = PRED7[20];
    PRED7_21_buffer[clk] = PRED7[21];
    PRED7_22_buffer[clk] = PRED7[22];
    PRED7_23_buffer[clk] = PRED7[23];
    PRED7_24_buffer[clk] = PRED7[24];
    PRED7_25_buffer[clk] = PRED7[25];
    PRED7_26_buffer[clk] = PRED7[26];
    PRED7_27_buffer[clk] = PRED7[27];
    PRED7_28_buffer[clk] = PRED7[28];
    PRED7_29_buffer[clk] = PRED7[29];
    PRED7_30_buffer[clk] = PRED7[30];
    PRED7_31_buffer[clk] = PRED7[31];
    PRED8_0_buffer[clk] = PRED8[0];
    PRED8_1_buffer[clk] = PRED8[1];
    PRED8_2_buffer[clk] = PRED8[2];
    PRED8_3_buffer[clk] = PRED8[3];
    PRED8_4_buffer[clk] = PRED8[4];
    PRED8_5_buffer[clk] = PRED8[5];
    PRED8_6_buffer[clk] = PRED8[6];
    PRED8_7_buffer[clk] = PRED8[7];
    PRED8_8_buffer[clk] = PRED8[8];
    PRED8_9_buffer[clk] = PRED8[9];
    PRED8_10_buffer[clk] = PRED8[10];
    PRED8_11_buffer[clk] = PRED8[11];
    PRED8_12_buffer[clk] = PRED8[12];
    PRED8_13_buffer[clk] = PRED8[13];
    PRED8_14_buffer[clk] = PRED8[14];
    PRED8_15_buffer[clk] = PRED8[15];
    PRED8_16_buffer[clk] = PRED8[16];
    PRED8_17_buffer[clk] = PRED8[17];
    PRED8_18_buffer[clk] = PRED8[18];
    PRED8_19_buffer[clk] = PRED8[19];
    PRED8_20_buffer[clk] = PRED8[20];
    PRED8_21_buffer[clk] = PRED8[21];
    PRED8_22_buffer[clk] = PRED8[22];
    PRED8_23_buffer[clk] = PRED8[23];
    PRED8_24_buffer[clk] = PRED8[24];
    PRED8_25_buffer[clk] = PRED8[25];
    PRED8_26_buffer[clk] = PRED8[26];
    PRED8_27_buffer[clk] = PRED8[27];
    PRED8_28_buffer[clk] = PRED8[28];
    PRED8_29_buffer[clk] = PRED8[29];
    PRED8_30_buffer[clk] = PRED8[30];
    PRED8_31_buffer[clk] = PRED8[31];
    PRED9_0_buffer[clk] = PRED9[0];
    PRED9_1_buffer[clk] = PRED9[1];
    PRED9_2_buffer[clk] = PRED9[2];
    PRED9_3_buffer[clk] = PRED9[3];
    PRED9_4_buffer[clk] = PRED9[4];
    PRED9_5_buffer[clk] = PRED9[5];
    PRED9_6_buffer[clk] = PRED9[6];
    PRED9_7_buffer[clk] = PRED9[7];
    PRED9_8_buffer[clk] = PRED9[8];
    PRED9_9_buffer[clk] = PRED9[9];
    PRED9_10_buffer[clk] = PRED9[10];
    PRED9_11_buffer[clk] = PRED9[11];
    PRED9_12_buffer[clk] = PRED9[12];
    PRED9_13_buffer[clk] = PRED9[13];
    PRED9_14_buffer[clk] = PRED9[14];
    PRED9_15_buffer[clk] = PRED9[15];
    PRED9_16_buffer[clk] = PRED9[16];
    PRED9_17_buffer[clk] = PRED9[17];
    PRED9_18_buffer[clk] = PRED9[18];
    PRED9_19_buffer[clk] = PRED9[19];
    PRED9_20_buffer[clk] = PRED9[20];
    PRED9_21_buffer[clk] = PRED9[21];
    PRED9_22_buffer[clk] = PRED9[22];
    PRED9_23_buffer[clk] = PRED9[23];
    PRED9_24_buffer[clk] = PRED9[24];
    PRED9_25_buffer[clk] = PRED9[25];
    PRED9_26_buffer[clk] = PRED9[26];
    PRED9_27_buffer[clk] = PRED9[27];
    PRED9_28_buffer[clk] = PRED9[28];
    PRED9_29_buffer[clk] = PRED9[29];
    PRED9_30_buffer[clk] = PRED9[30];
    PRED9_31_buffer[clk] = PRED9[31];
    PRED10_0_buffer[clk] = PRED10[0];
    PRED10_1_buffer[clk] = PRED10[1];
    PRED10_2_buffer[clk] = PRED10[2];
    PRED10_3_buffer[clk] = PRED10[3];
    PRED10_4_buffer[clk] = PRED10[4];
    PRED10_5_buffer[clk] = PRED10[5];
    PRED10_6_buffer[clk] = PRED10[6];
    PRED10_7_buffer[clk] = PRED10[7];
    PRED10_8_buffer[clk] = PRED10[8];
    PRED10_9_buffer[clk] = PRED10[9];
    PRED10_10_buffer[clk] = PRED10[10];
    PRED10_11_buffer[clk] = PRED10[11];
    PRED10_12_buffer[clk] = PRED10[12];
    PRED10_13_buffer[clk] = PRED10[13];
    PRED10_14_buffer[clk] = PRED10[14];
    PRED10_15_buffer[clk] = PRED10[15];
    PRED10_16_buffer[clk] = PRED10[16];
    PRED10_17_buffer[clk] = PRED10[17];
    PRED10_18_buffer[clk] = PRED10[18];
    PRED10_19_buffer[clk] = PRED10[19];
    PRED10_20_buffer[clk] = PRED10[20];
    PRED10_21_buffer[clk] = PRED10[21];
    PRED10_22_buffer[clk] = PRED10[22];
    PRED10_23_buffer[clk] = PRED10[23];
    PRED10_24_buffer[clk] = PRED10[24];
    PRED10_25_buffer[clk] = PRED10[25];
    PRED10_26_buffer[clk] = PRED10[26];
    PRED10_27_buffer[clk] = PRED10[27];
    PRED10_28_buffer[clk] = PRED10[28];
    PRED10_29_buffer[clk] = PRED10[29];
    PRED10_30_buffer[clk] = PRED10[30];
    PRED10_31_buffer[clk] = PRED10[31];
    PRED11_0_buffer[clk] = PRED11[0];
    PRED11_1_buffer[clk] = PRED11[1];
    PRED11_2_buffer[clk] = PRED11[2];
    PRED11_3_buffer[clk] = PRED11[3];
    PRED11_4_buffer[clk] = PRED11[4];
    PRED11_5_buffer[clk] = PRED11[5];
    PRED11_6_buffer[clk] = PRED11[6];
    PRED11_7_buffer[clk] = PRED11[7];
    PRED11_8_buffer[clk] = PRED11[8];
    PRED11_9_buffer[clk] = PRED11[9];
    PRED11_10_buffer[clk] = PRED11[10];
    PRED11_11_buffer[clk] = PRED11[11];
    PRED11_12_buffer[clk] = PRED11[12];
    PRED11_13_buffer[clk] = PRED11[13];
    PRED11_14_buffer[clk] = PRED11[14];
    PRED11_15_buffer[clk] = PRED11[15];
    PRED11_16_buffer[clk] = PRED11[16];
    PRED11_17_buffer[clk] = PRED11[17];
    PRED11_18_buffer[clk] = PRED11[18];
    PRED11_19_buffer[clk] = PRED11[19];
    PRED11_20_buffer[clk] = PRED11[20];
    PRED11_21_buffer[clk] = PRED11[21];
    PRED11_22_buffer[clk] = PRED11[22];
    PRED11_23_buffer[clk] = PRED11[23];
    PRED11_24_buffer[clk] = PRED11[24];
    PRED11_25_buffer[clk] = PRED11[25];
    PRED11_26_buffer[clk] = PRED11[26];
    PRED11_27_buffer[clk] = PRED11[27];
    PRED11_28_buffer[clk] = PRED11[28];
    PRED11_29_buffer[clk] = PRED11[29];
    PRED11_30_buffer[clk] = PRED11[30];
    PRED11_31_buffer[clk] = PRED11[31];
    PRED12_0_buffer[clk] = PRED12[0];
    PRED12_1_buffer[clk] = PRED12[1];
    PRED12_2_buffer[clk] = PRED12[2];
    PRED12_3_buffer[clk] = PRED12[3];
    PRED12_4_buffer[clk] = PRED12[4];
    PRED12_5_buffer[clk] = PRED12[5];
    PRED12_6_buffer[clk] = PRED12[6];
    PRED12_7_buffer[clk] = PRED12[7];
    PRED12_8_buffer[clk] = PRED12[8];
    PRED12_9_buffer[clk] = PRED12[9];
    PRED12_10_buffer[clk] = PRED12[10];
    PRED12_11_buffer[clk] = PRED12[11];
    PRED12_12_buffer[clk] = PRED12[12];
    PRED12_13_buffer[clk] = PRED12[13];
    PRED12_14_buffer[clk] = PRED12[14];
    PRED12_15_buffer[clk] = PRED12[15];
    PRED12_16_buffer[clk] = PRED12[16];
    PRED12_17_buffer[clk] = PRED12[17];
    PRED12_18_buffer[clk] = PRED12[18];
    PRED12_19_buffer[clk] = PRED12[19];
    PRED12_20_buffer[clk] = PRED12[20];
    PRED12_21_buffer[clk] = PRED12[21];
    PRED12_22_buffer[clk] = PRED12[22];
    PRED12_23_buffer[clk] = PRED12[23];
    PRED12_24_buffer[clk] = PRED12[24];
    PRED12_25_buffer[clk] = PRED12[25];
    PRED12_26_buffer[clk] = PRED12[26];
    PRED12_27_buffer[clk] = PRED12[27];
    PRED12_28_buffer[clk] = PRED12[28];
    PRED12_29_buffer[clk] = PRED12[29];
    PRED12_30_buffer[clk] = PRED12[30];
    PRED12_31_buffer[clk] = PRED12[31];
    PRED13_0_buffer[clk] = PRED13[0];
    PRED13_1_buffer[clk] = PRED13[1];
    PRED13_2_buffer[clk] = PRED13[2];
    PRED13_3_buffer[clk] = PRED13[3];
    PRED13_4_buffer[clk] = PRED13[4];
    PRED13_5_buffer[clk] = PRED13[5];
    PRED13_6_buffer[clk] = PRED13[6];
    PRED13_7_buffer[clk] = PRED13[7];
    PRED13_8_buffer[clk] = PRED13[8];
    PRED13_9_buffer[clk] = PRED13[9];
    PRED13_10_buffer[clk] = PRED13[10];
    PRED13_11_buffer[clk] = PRED13[11];
    PRED13_12_buffer[clk] = PRED13[12];
    PRED13_13_buffer[clk] = PRED13[13];
    PRED13_14_buffer[clk] = PRED13[14];
    PRED13_15_buffer[clk] = PRED13[15];
    PRED13_16_buffer[clk] = PRED13[16];
    PRED13_17_buffer[clk] = PRED13[17];
    PRED13_18_buffer[clk] = PRED13[18];
    PRED13_19_buffer[clk] = PRED13[19];
    PRED13_20_buffer[clk] = PRED13[20];
    PRED13_21_buffer[clk] = PRED13[21];
    PRED13_22_buffer[clk] = PRED13[22];
    PRED13_23_buffer[clk] = PRED13[23];
    PRED13_24_buffer[clk] = PRED13[24];
    PRED13_25_buffer[clk] = PRED13[25];
    PRED13_26_buffer[clk] = PRED13[26];
    PRED13_27_buffer[clk] = PRED13[27];
    PRED13_28_buffer[clk] = PRED13[28];
    PRED13_29_buffer[clk] = PRED13[29];
    PRED13_30_buffer[clk] = PRED13[30];
    PRED13_31_buffer[clk] = PRED13[31];
    PRED14_0_buffer[clk] = PRED14[0];
    PRED14_1_buffer[clk] = PRED14[1];
    PRED14_2_buffer[clk] = PRED14[2];
    PRED14_3_buffer[clk] = PRED14[3];
    PRED14_4_buffer[clk] = PRED14[4];
    PRED14_5_buffer[clk] = PRED14[5];
    PRED14_6_buffer[clk] = PRED14[6];
    PRED14_7_buffer[clk] = PRED14[7];
    PRED14_8_buffer[clk] = PRED14[8];
    PRED14_9_buffer[clk] = PRED14[9];
    PRED14_10_buffer[clk] = PRED14[10];
    PRED14_11_buffer[clk] = PRED14[11];
    PRED14_12_buffer[clk] = PRED14[12];
    PRED14_13_buffer[clk] = PRED14[13];
    PRED14_14_buffer[clk] = PRED14[14];
    PRED14_15_buffer[clk] = PRED14[15];
    PRED14_16_buffer[clk] = PRED14[16];
    PRED14_17_buffer[clk] = PRED14[17];
    PRED14_18_buffer[clk] = PRED14[18];
    PRED14_19_buffer[clk] = PRED14[19];
    PRED14_20_buffer[clk] = PRED14[20];
    PRED14_21_buffer[clk] = PRED14[21];
    PRED14_22_buffer[clk] = PRED14[22];
    PRED14_23_buffer[clk] = PRED14[23];
    PRED14_24_buffer[clk] = PRED14[24];
    PRED14_25_buffer[clk] = PRED14[25];
    PRED14_26_buffer[clk] = PRED14[26];
    PRED14_27_buffer[clk] = PRED14[27];
    PRED14_28_buffer[clk] = PRED14[28];
    PRED14_29_buffer[clk] = PRED14[29];
    PRED14_30_buffer[clk] = PRED14[30];
    PRED14_31_buffer[clk] = PRED14[31];
    PRED15_0_buffer[clk] = PRED15[0];
    PRED15_1_buffer[clk] = PRED15[1];
    PRED15_2_buffer[clk] = PRED15[2];
    PRED15_3_buffer[clk] = PRED15[3];
    PRED15_4_buffer[clk] = PRED15[4];
    PRED15_5_buffer[clk] = PRED15[5];
    PRED15_6_buffer[clk] = PRED15[6];
    PRED15_7_buffer[clk] = PRED15[7];
    PRED15_8_buffer[clk] = PRED15[8];
    PRED15_9_buffer[clk] = PRED15[9];
    PRED15_10_buffer[clk] = PRED15[10];
    PRED15_11_buffer[clk] = PRED15[11];
    PRED15_12_buffer[clk] = PRED15[12];
    PRED15_13_buffer[clk] = PRED15[13];
    PRED15_14_buffer[clk] = PRED15[14];
    PRED15_15_buffer[clk] = PRED15[15];
    PRED15_16_buffer[clk] = PRED15[16];
    PRED15_17_buffer[clk] = PRED15[17];
    PRED15_18_buffer[clk] = PRED15[18];
    PRED15_19_buffer[clk] = PRED15[19];
    PRED15_20_buffer[clk] = PRED15[20];
    PRED15_21_buffer[clk] = PRED15[21];
    PRED15_22_buffer[clk] = PRED15[22];
    PRED15_23_buffer[clk] = PRED15[23];
    PRED15_24_buffer[clk] = PRED15[24];
    PRED15_25_buffer[clk] = PRED15[25];
    PRED15_26_buffer[clk] = PRED15[26];
    PRED15_27_buffer[clk] = PRED15[27];
    PRED15_28_buffer[clk] = PRED15[28];
    PRED15_29_buffer[clk] = PRED15[29];
    PRED15_30_buffer[clk] = PRED15[30];
    PRED15_31_buffer[clk] = PRED15[31];
    PRED16_0_buffer[clk] = PRED16[0];
    PRED16_1_buffer[clk] = PRED16[1];
    PRED16_2_buffer[clk] = PRED16[2];
    PRED16_3_buffer[clk] = PRED16[3];
    PRED16_4_buffer[clk] = PRED16[4];
    PRED16_5_buffer[clk] = PRED16[5];
    PRED16_6_buffer[clk] = PRED16[6];
    PRED16_7_buffer[clk] = PRED16[7];
    PRED16_8_buffer[clk] = PRED16[8];
    PRED16_9_buffer[clk] = PRED16[9];
    PRED16_10_buffer[clk] = PRED16[10];
    PRED16_11_buffer[clk] = PRED16[11];
    PRED16_12_buffer[clk] = PRED16[12];
    PRED16_13_buffer[clk] = PRED16[13];
    PRED16_14_buffer[clk] = PRED16[14];
    PRED16_15_buffer[clk] = PRED16[15];
    PRED16_16_buffer[clk] = PRED16[16];
    PRED16_17_buffer[clk] = PRED16[17];
    PRED16_18_buffer[clk] = PRED16[18];
    PRED16_19_buffer[clk] = PRED16[19];
    PRED16_20_buffer[clk] = PRED16[20];
    PRED16_21_buffer[clk] = PRED16[21];
    PRED16_22_buffer[clk] = PRED16[22];
    PRED16_23_buffer[clk] = PRED16[23];
    PRED16_24_buffer[clk] = PRED16[24];
    PRED16_25_buffer[clk] = PRED16[25];
    PRED16_26_buffer[clk] = PRED16[26];
    PRED16_27_buffer[clk] = PRED16[27];
    PRED16_28_buffer[clk] = PRED16[28];
    PRED16_29_buffer[clk] = PRED16[29];
    PRED16_30_buffer[clk] = PRED16[30];
    PRED16_31_buffer[clk] = PRED16[31];
    PRED17_0_buffer[clk] = PRED17[0];
    PRED17_1_buffer[clk] = PRED17[1];
    PRED17_2_buffer[clk] = PRED17[2];
    PRED17_3_buffer[clk] = PRED17[3];
    PRED17_4_buffer[clk] = PRED17[4];
    PRED17_5_buffer[clk] = PRED17[5];
    PRED17_6_buffer[clk] = PRED17[6];
    PRED17_7_buffer[clk] = PRED17[7];
    PRED17_8_buffer[clk] = PRED17[8];
    PRED17_9_buffer[clk] = PRED17[9];
    PRED17_10_buffer[clk] = PRED17[10];
    PRED17_11_buffer[clk] = PRED17[11];
    PRED17_12_buffer[clk] = PRED17[12];
    PRED17_13_buffer[clk] = PRED17[13];
    PRED17_14_buffer[clk] = PRED17[14];
    PRED17_15_buffer[clk] = PRED17[15];
    PRED17_16_buffer[clk] = PRED17[16];
    PRED17_17_buffer[clk] = PRED17[17];
    PRED17_18_buffer[clk] = PRED17[18];
    PRED17_19_buffer[clk] = PRED17[19];
    PRED17_20_buffer[clk] = PRED17[20];
    PRED17_21_buffer[clk] = PRED17[21];
    PRED17_22_buffer[clk] = PRED17[22];
    PRED17_23_buffer[clk] = PRED17[23];
    PRED17_24_buffer[clk] = PRED17[24];
    PRED17_25_buffer[clk] = PRED17[25];
    PRED17_26_buffer[clk] = PRED17[26];
    PRED17_27_buffer[clk] = PRED17[27];
    PRED17_28_buffer[clk] = PRED17[28];
    PRED17_29_buffer[clk] = PRED17[29];
    PRED17_30_buffer[clk] = PRED17[30];
    PRED17_31_buffer[clk] = PRED17[31];
    PRED18_0_buffer[clk] = PRED18[0];
    PRED18_1_buffer[clk] = PRED18[1];
    PRED18_2_buffer[clk] = PRED18[2];
    PRED18_3_buffer[clk] = PRED18[3];
    PRED18_4_buffer[clk] = PRED18[4];
    PRED18_5_buffer[clk] = PRED18[5];
    PRED18_6_buffer[clk] = PRED18[6];
    PRED18_7_buffer[clk] = PRED18[7];
    PRED18_8_buffer[clk] = PRED18[8];
    PRED18_9_buffer[clk] = PRED18[9];
    PRED18_10_buffer[clk] = PRED18[10];
    PRED18_11_buffer[clk] = PRED18[11];
    PRED18_12_buffer[clk] = PRED18[12];
    PRED18_13_buffer[clk] = PRED18[13];
    PRED18_14_buffer[clk] = PRED18[14];
    PRED18_15_buffer[clk] = PRED18[15];
    PRED18_16_buffer[clk] = PRED18[16];
    PRED18_17_buffer[clk] = PRED18[17];
    PRED18_18_buffer[clk] = PRED18[18];
    PRED18_19_buffer[clk] = PRED18[19];
    PRED18_20_buffer[clk] = PRED18[20];
    PRED18_21_buffer[clk] = PRED18[21];
    PRED18_22_buffer[clk] = PRED18[22];
    PRED18_23_buffer[clk] = PRED18[23];
    PRED18_24_buffer[clk] = PRED18[24];
    PRED18_25_buffer[clk] = PRED18[25];
    PRED18_26_buffer[clk] = PRED18[26];
    PRED18_27_buffer[clk] = PRED18[27];
    PRED18_28_buffer[clk] = PRED18[28];
    PRED18_29_buffer[clk] = PRED18[29];
    PRED18_30_buffer[clk] = PRED18[30];
    PRED18_31_buffer[clk] = PRED18[31];
    PRED19_0_buffer[clk] = PRED19[0];
    PRED19_1_buffer[clk] = PRED19[1];
    PRED19_2_buffer[clk] = PRED19[2];
    PRED19_3_buffer[clk] = PRED19[3];
    PRED19_4_buffer[clk] = PRED19[4];
    PRED19_5_buffer[clk] = PRED19[5];
    PRED19_6_buffer[clk] = PRED19[6];
    PRED19_7_buffer[clk] = PRED19[7];
    PRED19_8_buffer[clk] = PRED19[8];
    PRED19_9_buffer[clk] = PRED19[9];
    PRED19_10_buffer[clk] = PRED19[10];
    PRED19_11_buffer[clk] = PRED19[11];
    PRED19_12_buffer[clk] = PRED19[12];
    PRED19_13_buffer[clk] = PRED19[13];
    PRED19_14_buffer[clk] = PRED19[14];
    PRED19_15_buffer[clk] = PRED19[15];
    PRED19_16_buffer[clk] = PRED19[16];
    PRED19_17_buffer[clk] = PRED19[17];
    PRED19_18_buffer[clk] = PRED19[18];
    PRED19_19_buffer[clk] = PRED19[19];
    PRED19_20_buffer[clk] = PRED19[20];
    PRED19_21_buffer[clk] = PRED19[21];
    PRED19_22_buffer[clk] = PRED19[22];
    PRED19_23_buffer[clk] = PRED19[23];
    PRED19_24_buffer[clk] = PRED19[24];
    PRED19_25_buffer[clk] = PRED19[25];
    PRED19_26_buffer[clk] = PRED19[26];
    PRED19_27_buffer[clk] = PRED19[27];
    PRED19_28_buffer[clk] = PRED19[28];
    PRED19_29_buffer[clk] = PRED19[29];
    PRED19_30_buffer[clk] = PRED19[30];
    PRED19_31_buffer[clk] = PRED19[31];
    PRED20_0_buffer[clk] = PRED20[0];
    PRED20_1_buffer[clk] = PRED20[1];
    PRED20_2_buffer[clk] = PRED20[2];
    PRED20_3_buffer[clk] = PRED20[3];
    PRED20_4_buffer[clk] = PRED20[4];
    PRED20_5_buffer[clk] = PRED20[5];
    PRED20_6_buffer[clk] = PRED20[6];
    PRED20_7_buffer[clk] = PRED20[7];
    PRED20_8_buffer[clk] = PRED20[8];
    PRED20_9_buffer[clk] = PRED20[9];
    PRED20_10_buffer[clk] = PRED20[10];
    PRED20_11_buffer[clk] = PRED20[11];
    PRED20_12_buffer[clk] = PRED20[12];
    PRED20_13_buffer[clk] = PRED20[13];
    PRED20_14_buffer[clk] = PRED20[14];
    PRED20_15_buffer[clk] = PRED20[15];
    PRED20_16_buffer[clk] = PRED20[16];
    PRED20_17_buffer[clk] = PRED20[17];
    PRED20_18_buffer[clk] = PRED20[18];
    PRED20_19_buffer[clk] = PRED20[19];
    PRED20_20_buffer[clk] = PRED20[20];
    PRED20_21_buffer[clk] = PRED20[21];
    PRED20_22_buffer[clk] = PRED20[22];
    PRED20_23_buffer[clk] = PRED20[23];
    PRED20_24_buffer[clk] = PRED20[24];
    PRED20_25_buffer[clk] = PRED20[25];
    PRED20_26_buffer[clk] = PRED20[26];
    PRED20_27_buffer[clk] = PRED20[27];
    PRED20_28_buffer[clk] = PRED20[28];
    PRED20_29_buffer[clk] = PRED20[29];
    PRED20_30_buffer[clk] = PRED20[30];
    PRED20_31_buffer[clk] = PRED20[31];
    PRED21_0_buffer[clk] = PRED21[0];
    PRED21_1_buffer[clk] = PRED21[1];
    PRED21_2_buffer[clk] = PRED21[2];
    PRED21_3_buffer[clk] = PRED21[3];
    PRED21_4_buffer[clk] = PRED21[4];
    PRED21_5_buffer[clk] = PRED21[5];
    PRED21_6_buffer[clk] = PRED21[6];
    PRED21_7_buffer[clk] = PRED21[7];
    PRED21_8_buffer[clk] = PRED21[8];
    PRED21_9_buffer[clk] = PRED21[9];
    PRED21_10_buffer[clk] = PRED21[10];
    PRED21_11_buffer[clk] = PRED21[11];
    PRED21_12_buffer[clk] = PRED21[12];
    PRED21_13_buffer[clk] = PRED21[13];
    PRED21_14_buffer[clk] = PRED21[14];
    PRED21_15_buffer[clk] = PRED21[15];
    PRED21_16_buffer[clk] = PRED21[16];
    PRED21_17_buffer[clk] = PRED21[17];
    PRED21_18_buffer[clk] = PRED21[18];
    PRED21_19_buffer[clk] = PRED21[19];
    PRED21_20_buffer[clk] = PRED21[20];
    PRED21_21_buffer[clk] = PRED21[21];
    PRED21_22_buffer[clk] = PRED21[22];
    PRED21_23_buffer[clk] = PRED21[23];
    PRED21_24_buffer[clk] = PRED21[24];
    PRED21_25_buffer[clk] = PRED21[25];
    PRED21_26_buffer[clk] = PRED21[26];
    PRED21_27_buffer[clk] = PRED21[27];
    PRED21_28_buffer[clk] = PRED21[28];
    PRED21_29_buffer[clk] = PRED21[29];
    PRED21_30_buffer[clk] = PRED21[30];
    PRED21_31_buffer[clk] = PRED21[31];
    PRED22_0_buffer[clk] = PRED22[0];
    PRED22_1_buffer[clk] = PRED22[1];
    PRED22_2_buffer[clk] = PRED22[2];
    PRED22_3_buffer[clk] = PRED22[3];
    PRED22_4_buffer[clk] = PRED22[4];
    PRED22_5_buffer[clk] = PRED22[5];
    PRED22_6_buffer[clk] = PRED22[6];
    PRED22_7_buffer[clk] = PRED22[7];
    PRED22_8_buffer[clk] = PRED22[8];
    PRED22_9_buffer[clk] = PRED22[9];
    PRED22_10_buffer[clk] = PRED22[10];
    PRED22_11_buffer[clk] = PRED22[11];
    PRED22_12_buffer[clk] = PRED22[12];
    PRED22_13_buffer[clk] = PRED22[13];
    PRED22_14_buffer[clk] = PRED22[14];
    PRED22_15_buffer[clk] = PRED22[15];
    PRED22_16_buffer[clk] = PRED22[16];
    PRED22_17_buffer[clk] = PRED22[17];
    PRED22_18_buffer[clk] = PRED22[18];
    PRED22_19_buffer[clk] = PRED22[19];
    PRED22_20_buffer[clk] = PRED22[20];
    PRED22_21_buffer[clk] = PRED22[21];
    PRED22_22_buffer[clk] = PRED22[22];
    PRED22_23_buffer[clk] = PRED22[23];
    PRED22_24_buffer[clk] = PRED22[24];
    PRED22_25_buffer[clk] = PRED22[25];
    PRED22_26_buffer[clk] = PRED22[26];
    PRED22_27_buffer[clk] = PRED22[27];
    PRED22_28_buffer[clk] = PRED22[28];
    PRED22_29_buffer[clk] = PRED22[29];
    PRED22_30_buffer[clk] = PRED22[30];
    PRED22_31_buffer[clk] = PRED22[31];
    PRED23_0_buffer[clk] = PRED23[0];
    PRED23_1_buffer[clk] = PRED23[1];
    PRED23_2_buffer[clk] = PRED23[2];
    PRED23_3_buffer[clk] = PRED23[3];
    PRED23_4_buffer[clk] = PRED23[4];
    PRED23_5_buffer[clk] = PRED23[5];
    PRED23_6_buffer[clk] = PRED23[6];
    PRED23_7_buffer[clk] = PRED23[7];
    PRED23_8_buffer[clk] = PRED23[8];
    PRED23_9_buffer[clk] = PRED23[9];
    PRED23_10_buffer[clk] = PRED23[10];
    PRED23_11_buffer[clk] = PRED23[11];
    PRED23_12_buffer[clk] = PRED23[12];
    PRED23_13_buffer[clk] = PRED23[13];
    PRED23_14_buffer[clk] = PRED23[14];
    PRED23_15_buffer[clk] = PRED23[15];
    PRED23_16_buffer[clk] = PRED23[16];
    PRED23_17_buffer[clk] = PRED23[17];
    PRED23_18_buffer[clk] = PRED23[18];
    PRED23_19_buffer[clk] = PRED23[19];
    PRED23_20_buffer[clk] = PRED23[20];
    PRED23_21_buffer[clk] = PRED23[21];
    PRED23_22_buffer[clk] = PRED23[22];
    PRED23_23_buffer[clk] = PRED23[23];
    PRED23_24_buffer[clk] = PRED23[24];
    PRED23_25_buffer[clk] = PRED23[25];
    PRED23_26_buffer[clk] = PRED23[26];
    PRED23_27_buffer[clk] = PRED23[27];
    PRED23_28_buffer[clk] = PRED23[28];
    PRED23_29_buffer[clk] = PRED23[29];
    PRED23_30_buffer[clk] = PRED23[30];
    PRED23_31_buffer[clk] = PRED23[31];
    PRED24_0_buffer[clk] = PRED24[0];
    PRED24_1_buffer[clk] = PRED24[1];
    PRED24_2_buffer[clk] = PRED24[2];
    PRED24_3_buffer[clk] = PRED24[3];
    PRED24_4_buffer[clk] = PRED24[4];
    PRED24_5_buffer[clk] = PRED24[5];
    PRED24_6_buffer[clk] = PRED24[6];
    PRED24_7_buffer[clk] = PRED24[7];
    PRED24_8_buffer[clk] = PRED24[8];
    PRED24_9_buffer[clk] = PRED24[9];
    PRED24_10_buffer[clk] = PRED24[10];
    PRED24_11_buffer[clk] = PRED24[11];
    PRED24_12_buffer[clk] = PRED24[12];
    PRED24_13_buffer[clk] = PRED24[13];
    PRED24_14_buffer[clk] = PRED24[14];
    PRED24_15_buffer[clk] = PRED24[15];
    PRED24_16_buffer[clk] = PRED24[16];
    PRED24_17_buffer[clk] = PRED24[17];
    PRED24_18_buffer[clk] = PRED24[18];
    PRED24_19_buffer[clk] = PRED24[19];
    PRED24_20_buffer[clk] = PRED24[20];
    PRED24_21_buffer[clk] = PRED24[21];
    PRED24_22_buffer[clk] = PRED24[22];
    PRED24_23_buffer[clk] = PRED24[23];
    PRED24_24_buffer[clk] = PRED24[24];
    PRED24_25_buffer[clk] = PRED24[25];
    PRED24_26_buffer[clk] = PRED24[26];
    PRED24_27_buffer[clk] = PRED24[27];
    PRED24_28_buffer[clk] = PRED24[28];
    PRED24_29_buffer[clk] = PRED24[29];
    PRED24_30_buffer[clk] = PRED24[30];
    PRED24_31_buffer[clk] = PRED24[31];
    PRED25_0_buffer[clk] = PRED25[0];
    PRED25_1_buffer[clk] = PRED25[1];
    PRED25_2_buffer[clk] = PRED25[2];
    PRED25_3_buffer[clk] = PRED25[3];
    PRED25_4_buffer[clk] = PRED25[4];
    PRED25_5_buffer[clk] = PRED25[5];
    PRED25_6_buffer[clk] = PRED25[6];
    PRED25_7_buffer[clk] = PRED25[7];
    PRED25_8_buffer[clk] = PRED25[8];
    PRED25_9_buffer[clk] = PRED25[9];
    PRED25_10_buffer[clk] = PRED25[10];
    PRED25_11_buffer[clk] = PRED25[11];
    PRED25_12_buffer[clk] = PRED25[12];
    PRED25_13_buffer[clk] = PRED25[13];
    PRED25_14_buffer[clk] = PRED25[14];
    PRED25_15_buffer[clk] = PRED25[15];
    PRED25_16_buffer[clk] = PRED25[16];
    PRED25_17_buffer[clk] = PRED25[17];
    PRED25_18_buffer[clk] = PRED25[18];
    PRED25_19_buffer[clk] = PRED25[19];
    PRED25_20_buffer[clk] = PRED25[20];
    PRED25_21_buffer[clk] = PRED25[21];
    PRED25_22_buffer[clk] = PRED25[22];
    PRED25_23_buffer[clk] = PRED25[23];
    PRED25_24_buffer[clk] = PRED25[24];
    PRED25_25_buffer[clk] = PRED25[25];
    PRED25_26_buffer[clk] = PRED25[26];
    PRED25_27_buffer[clk] = PRED25[27];
    PRED25_28_buffer[clk] = PRED25[28];
    PRED25_29_buffer[clk] = PRED25[29];
    PRED25_30_buffer[clk] = PRED25[30];
    PRED25_31_buffer[clk] = PRED25[31];
    PRED26_0_buffer[clk] = PRED26[0];
    PRED26_1_buffer[clk] = PRED26[1];
    PRED26_2_buffer[clk] = PRED26[2];
    PRED26_3_buffer[clk] = PRED26[3];
    PRED26_4_buffer[clk] = PRED26[4];
    PRED26_5_buffer[clk] = PRED26[5];
    PRED26_6_buffer[clk] = PRED26[6];
    PRED26_7_buffer[clk] = PRED26[7];
    PRED26_8_buffer[clk] = PRED26[8];
    PRED26_9_buffer[clk] = PRED26[9];
    PRED26_10_buffer[clk] = PRED26[10];
    PRED26_11_buffer[clk] = PRED26[11];
    PRED26_12_buffer[clk] = PRED26[12];
    PRED26_13_buffer[clk] = PRED26[13];
    PRED26_14_buffer[clk] = PRED26[14];
    PRED26_15_buffer[clk] = PRED26[15];
    PRED26_16_buffer[clk] = PRED26[16];
    PRED26_17_buffer[clk] = PRED26[17];
    PRED26_18_buffer[clk] = PRED26[18];
    PRED26_19_buffer[clk] = PRED26[19];
    PRED26_20_buffer[clk] = PRED26[20];
    PRED26_21_buffer[clk] = PRED26[21];
    PRED26_22_buffer[clk] = PRED26[22];
    PRED26_23_buffer[clk] = PRED26[23];
    PRED26_24_buffer[clk] = PRED26[24];
    PRED26_25_buffer[clk] = PRED26[25];
    PRED26_26_buffer[clk] = PRED26[26];
    PRED26_27_buffer[clk] = PRED26[27];
    PRED26_28_buffer[clk] = PRED26[28];
    PRED26_29_buffer[clk] = PRED26[29];
    PRED26_30_buffer[clk] = PRED26[30];
    PRED26_31_buffer[clk] = PRED26[31];
    PRED27_0_buffer[clk] = PRED27[0];
    PRED27_1_buffer[clk] = PRED27[1];
    PRED27_2_buffer[clk] = PRED27[2];
    PRED27_3_buffer[clk] = PRED27[3];
    PRED27_4_buffer[clk] = PRED27[4];
    PRED27_5_buffer[clk] = PRED27[5];
    PRED27_6_buffer[clk] = PRED27[6];
    PRED27_7_buffer[clk] = PRED27[7];
    PRED27_8_buffer[clk] = PRED27[8];
    PRED27_9_buffer[clk] = PRED27[9];
    PRED27_10_buffer[clk] = PRED27[10];
    PRED27_11_buffer[clk] = PRED27[11];
    PRED27_12_buffer[clk] = PRED27[12];
    PRED27_13_buffer[clk] = PRED27[13];
    PRED27_14_buffer[clk] = PRED27[14];
    PRED27_15_buffer[clk] = PRED27[15];
    PRED27_16_buffer[clk] = PRED27[16];
    PRED27_17_buffer[clk] = PRED27[17];
    PRED27_18_buffer[clk] = PRED27[18];
    PRED27_19_buffer[clk] = PRED27[19];
    PRED27_20_buffer[clk] = PRED27[20];
    PRED27_21_buffer[clk] = PRED27[21];
    PRED27_22_buffer[clk] = PRED27[22];
    PRED27_23_buffer[clk] = PRED27[23];
    PRED27_24_buffer[clk] = PRED27[24];
    PRED27_25_buffer[clk] = PRED27[25];
    PRED27_26_buffer[clk] = PRED27[26];
    PRED27_27_buffer[clk] = PRED27[27];
    PRED27_28_buffer[clk] = PRED27[28];
    PRED27_29_buffer[clk] = PRED27[29];
    PRED27_30_buffer[clk] = PRED27[30];
    PRED27_31_buffer[clk] = PRED27[31];
    PRED28_0_buffer[clk] = PRED28[0];
    PRED28_1_buffer[clk] = PRED28[1];
    PRED28_2_buffer[clk] = PRED28[2];
    PRED28_3_buffer[clk] = PRED28[3];
    PRED28_4_buffer[clk] = PRED28[4];
    PRED28_5_buffer[clk] = PRED28[5];
    PRED28_6_buffer[clk] = PRED28[6];
    PRED28_7_buffer[clk] = PRED28[7];
    PRED28_8_buffer[clk] = PRED28[8];
    PRED28_9_buffer[clk] = PRED28[9];
    PRED28_10_buffer[clk] = PRED28[10];
    PRED28_11_buffer[clk] = PRED28[11];
    PRED28_12_buffer[clk] = PRED28[12];
    PRED28_13_buffer[clk] = PRED28[13];
    PRED28_14_buffer[clk] = PRED28[14];
    PRED28_15_buffer[clk] = PRED28[15];
    PRED28_16_buffer[clk] = PRED28[16];
    PRED28_17_buffer[clk] = PRED28[17];
    PRED28_18_buffer[clk] = PRED28[18];
    PRED28_19_buffer[clk] = PRED28[19];
    PRED28_20_buffer[clk] = PRED28[20];
    PRED28_21_buffer[clk] = PRED28[21];
    PRED28_22_buffer[clk] = PRED28[22];
    PRED28_23_buffer[clk] = PRED28[23];
    PRED28_24_buffer[clk] = PRED28[24];
    PRED28_25_buffer[clk] = PRED28[25];
    PRED28_26_buffer[clk] = PRED28[26];
    PRED28_27_buffer[clk] = PRED28[27];
    PRED28_28_buffer[clk] = PRED28[28];
    PRED28_29_buffer[clk] = PRED28[29];
    PRED28_30_buffer[clk] = PRED28[30];
    PRED28_31_buffer[clk] = PRED28[31];
    PRED29_0_buffer[clk] = PRED29[0];
    PRED29_1_buffer[clk] = PRED29[1];
    PRED29_2_buffer[clk] = PRED29[2];
    PRED29_3_buffer[clk] = PRED29[3];
    PRED29_4_buffer[clk] = PRED29[4];
    PRED29_5_buffer[clk] = PRED29[5];
    PRED29_6_buffer[clk] = PRED29[6];
    PRED29_7_buffer[clk] = PRED29[7];
    PRED29_8_buffer[clk] = PRED29[8];
    PRED29_9_buffer[clk] = PRED29[9];
    PRED29_10_buffer[clk] = PRED29[10];
    PRED29_11_buffer[clk] = PRED29[11];
    PRED29_12_buffer[clk] = PRED29[12];
    PRED29_13_buffer[clk] = PRED29[13];
    PRED29_14_buffer[clk] = PRED29[14];
    PRED29_15_buffer[clk] = PRED29[15];
    PRED29_16_buffer[clk] = PRED29[16];
    PRED29_17_buffer[clk] = PRED29[17];
    PRED29_18_buffer[clk] = PRED29[18];
    PRED29_19_buffer[clk] = PRED29[19];
    PRED29_20_buffer[clk] = PRED29[20];
    PRED29_21_buffer[clk] = PRED29[21];
    PRED29_22_buffer[clk] = PRED29[22];
    PRED29_23_buffer[clk] = PRED29[23];
    PRED29_24_buffer[clk] = PRED29[24];
    PRED29_25_buffer[clk] = PRED29[25];
    PRED29_26_buffer[clk] = PRED29[26];
    PRED29_27_buffer[clk] = PRED29[27];
    PRED29_28_buffer[clk] = PRED29[28];
    PRED29_29_buffer[clk] = PRED29[29];
    PRED29_30_buffer[clk] = PRED29[30];
    PRED29_31_buffer[clk] = PRED29[31];
    PRED30_0_buffer[clk] = PRED30[0];
    PRED30_1_buffer[clk] = PRED30[1];
    PRED30_2_buffer[clk] = PRED30[2];
    PRED30_3_buffer[clk] = PRED30[3];
    PRED30_4_buffer[clk] = PRED30[4];
    PRED30_5_buffer[clk] = PRED30[5];
    PRED30_6_buffer[clk] = PRED30[6];
    PRED30_7_buffer[clk] = PRED30[7];
    PRED30_8_buffer[clk] = PRED30[8];
    PRED30_9_buffer[clk] = PRED30[9];
    PRED30_10_buffer[clk] = PRED30[10];
    PRED30_11_buffer[clk] = PRED30[11];
    PRED30_12_buffer[clk] = PRED30[12];
    PRED30_13_buffer[clk] = PRED30[13];
    PRED30_14_buffer[clk] = PRED30[14];
    PRED30_15_buffer[clk] = PRED30[15];
    PRED30_16_buffer[clk] = PRED30[16];
    PRED30_17_buffer[clk] = PRED30[17];
    PRED30_18_buffer[clk] = PRED30[18];
    PRED30_19_buffer[clk] = PRED30[19];
    PRED30_20_buffer[clk] = PRED30[20];
    PRED30_21_buffer[clk] = PRED30[21];
    PRED30_22_buffer[clk] = PRED30[22];
    PRED30_23_buffer[clk] = PRED30[23];
    PRED30_24_buffer[clk] = PRED30[24];
    PRED30_25_buffer[clk] = PRED30[25];
    PRED30_26_buffer[clk] = PRED30[26];
    PRED30_27_buffer[clk] = PRED30[27];
    PRED30_28_buffer[clk] = PRED30[28];
    PRED30_29_buffer[clk] = PRED30[29];
    PRED30_30_buffer[clk] = PRED30[30];
    PRED30_31_buffer[clk] = PRED30[31];
    PRED31_0_buffer[clk] = PRED31[0];
    PRED31_1_buffer[clk] = PRED31[1];
    PRED31_2_buffer[clk] = PRED31[2];
    PRED31_3_buffer[clk] = PRED31[3];
    PRED31_4_buffer[clk] = PRED31[4];
    PRED31_5_buffer[clk] = PRED31[5];
    PRED31_6_buffer[clk] = PRED31[6];
    PRED31_7_buffer[clk] = PRED31[7];
    PRED31_8_buffer[clk] = PRED31[8];
    PRED31_9_buffer[clk] = PRED31[9];
    PRED31_10_buffer[clk] = PRED31[10];
    PRED31_11_buffer[clk] = PRED31[11];
    PRED31_12_buffer[clk] = PRED31[12];
    PRED31_13_buffer[clk] = PRED31[13];
    PRED31_14_buffer[clk] = PRED31[14];
    PRED31_15_buffer[clk] = PRED31[15];
    PRED31_16_buffer[clk] = PRED31[16];
    PRED31_17_buffer[clk] = PRED31[17];
    PRED31_18_buffer[clk] = PRED31[18];
    PRED31_19_buffer[clk] = PRED31[19];
    PRED31_20_buffer[clk] = PRED31[20];
    PRED31_21_buffer[clk] = PRED31[21];
    PRED31_22_buffer[clk] = PRED31[22];
    PRED31_23_buffer[clk] = PRED31[23];
    PRED31_24_buffer[clk] = PRED31[24];
    PRED31_25_buffer[clk] = PRED31[25];
    PRED31_26_buffer[clk] = PRED31[26];
    PRED31_27_buffer[clk] = PRED31[27];
    PRED31_28_buffer[clk] = PRED31[28];
    PRED31_29_buffer[clk] = PRED31[29];
    PRED31_30_buffer[clk] = PRED31[30];
    PRED31_31_buffer[clk] = PRED31[31];
    PRED32_0_buffer[clk] = PRED32[0];
    PRED32_1_buffer[clk] = PRED32[1];
    PRED32_2_buffer[clk] = PRED32[2];
    PRED32_3_buffer[clk] = PRED32[3];
    PRED32_4_buffer[clk] = PRED32[4];
    PRED32_5_buffer[clk] = PRED32[5];
    PRED32_6_buffer[clk] = PRED32[6];
    PRED32_7_buffer[clk] = PRED32[7];
    PRED32_8_buffer[clk] = PRED32[8];
    PRED32_9_buffer[clk] = PRED32[9];
    PRED32_10_buffer[clk] = PRED32[10];
    PRED32_11_buffer[clk] = PRED32[11];
    PRED32_12_buffer[clk] = PRED32[12];
    PRED32_13_buffer[clk] = PRED32[13];
    PRED32_14_buffer[clk] = PRED32[14];
    PRED32_15_buffer[clk] = PRED32[15];
    PRED32_16_buffer[clk] = PRED32[16];
    PRED32_17_buffer[clk] = PRED32[17];
    PRED32_18_buffer[clk] = PRED32[18];
    PRED32_19_buffer[clk] = PRED32[19];
    PRED32_20_buffer[clk] = PRED32[20];
    PRED32_21_buffer[clk] = PRED32[21];
    PRED32_22_buffer[clk] = PRED32[22];
    PRED32_23_buffer[clk] = PRED32[23];
    PRED32_24_buffer[clk] = PRED32[24];
    PRED32_25_buffer[clk] = PRED32[25];
    PRED32_26_buffer[clk] = PRED32[26];
    PRED32_27_buffer[clk] = PRED32[27];
    PRED32_28_buffer[clk] = PRED32[28];
    PRED32_29_buffer[clk] = PRED32[29];
    PRED32_30_buffer[clk] = PRED32[30];
    PRED32_31_buffer[clk] = PRED32[31];
    PRED33_0_buffer[clk] = PRED33[0];
    PRED33_1_buffer[clk] = PRED33[1];
    PRED33_2_buffer[clk] = PRED33[2];
    PRED33_3_buffer[clk] = PRED33[3];
    PRED33_4_buffer[clk] = PRED33[4];
    PRED33_5_buffer[clk] = PRED33[5];
    PRED33_6_buffer[clk] = PRED33[6];
    PRED33_7_buffer[clk] = PRED33[7];
    PRED33_8_buffer[clk] = PRED33[8];
    PRED33_9_buffer[clk] = PRED33[9];
    PRED33_10_buffer[clk] = PRED33[10];
    PRED33_11_buffer[clk] = PRED33[11];
    PRED33_12_buffer[clk] = PRED33[12];
    PRED33_13_buffer[clk] = PRED33[13];
    PRED33_14_buffer[clk] = PRED33[14];
    PRED33_15_buffer[clk] = PRED33[15];
    PRED33_16_buffer[clk] = PRED33[16];
    PRED33_17_buffer[clk] = PRED33[17];
    PRED33_18_buffer[clk] = PRED33[18];
    PRED33_19_buffer[clk] = PRED33[19];
    PRED33_20_buffer[clk] = PRED33[20];
    PRED33_21_buffer[clk] = PRED33[21];
    PRED33_22_buffer[clk] = PRED33[22];
    PRED33_23_buffer[clk] = PRED33[23];
    PRED33_24_buffer[clk] = PRED33[24];
    PRED33_25_buffer[clk] = PRED33[25];
    PRED33_26_buffer[clk] = PRED33[26];
    PRED33_27_buffer[clk] = PRED33[27];
    PRED33_28_buffer[clk] = PRED33[28];
    PRED33_29_buffer[clk] = PRED33[29];
    PRED33_30_buffer[clk] = PRED33[30];
    PRED33_31_buffer[clk] = PRED33[31];
    PRED34_0_buffer[clk] = PRED34[0];
    PRED34_1_buffer[clk] = PRED34[1];
    PRED34_2_buffer[clk] = PRED34[2];
    PRED34_3_buffer[clk] = PRED34[3];
    PRED34_4_buffer[clk] = PRED34[4];
    PRED34_5_buffer[clk] = PRED34[5];
    PRED34_6_buffer[clk] = PRED34[6];
    PRED34_7_buffer[clk] = PRED34[7];
    PRED34_8_buffer[clk] = PRED34[8];
    PRED34_9_buffer[clk] = PRED34[9];
    PRED34_10_buffer[clk] = PRED34[10];
    PRED34_11_buffer[clk] = PRED34[11];
    PRED34_12_buffer[clk] = PRED34[12];
    PRED34_13_buffer[clk] = PRED34[13];
    PRED34_14_buffer[clk] = PRED34[14];
    PRED34_15_buffer[clk] = PRED34[15];
    PRED34_16_buffer[clk] = PRED34[16];
    PRED34_17_buffer[clk] = PRED34[17];
    PRED34_18_buffer[clk] = PRED34[18];
    PRED34_19_buffer[clk] = PRED34[19];
    PRED34_20_buffer[clk] = PRED34[20];
    PRED34_21_buffer[clk] = PRED34[21];
    PRED34_22_buffer[clk] = PRED34[22];
    PRED34_23_buffer[clk] = PRED34[23];
    PRED34_24_buffer[clk] = PRED34[24];
    PRED34_25_buffer[clk] = PRED34[25];
    PRED34_26_buffer[clk] = PRED34[26];
    PRED34_27_buffer[clk] = PRED34[27];
    PRED34_28_buffer[clk] = PRED34[28];
    PRED34_29_buffer[clk] = PRED34[29];
    PRED34_30_buffer[clk] = PRED34[30];
    PRED34_31_buffer[clk] = PRED34[31];
    PRED35_0_buffer[clk] = PRED35[0];
    PRED35_1_buffer[clk] = PRED35[1];
    PRED35_2_buffer[clk] = PRED35[2];
    PRED35_3_buffer[clk] = PRED35[3];
    PRED35_4_buffer[clk] = PRED35[4];
    PRED35_5_buffer[clk] = PRED35[5];
    PRED35_6_buffer[clk] = PRED35[6];
    PRED35_7_buffer[clk] = PRED35[7];
    PRED35_8_buffer[clk] = PRED35[8];
    PRED35_9_buffer[clk] = PRED35[9];
    PRED35_10_buffer[clk] = PRED35[10];
    PRED35_11_buffer[clk] = PRED35[11];
    PRED35_12_buffer[clk] = PRED35[12];
    PRED35_13_buffer[clk] = PRED35[13];
    PRED35_14_buffer[clk] = PRED35[14];
    PRED35_15_buffer[clk] = PRED35[15];
    PRED35_16_buffer[clk] = PRED35[16];
    PRED35_17_buffer[clk] = PRED35[17];
    PRED35_18_buffer[clk] = PRED35[18];
    PRED35_19_buffer[clk] = PRED35[19];
    PRED35_20_buffer[clk] = PRED35[20];
    PRED35_21_buffer[clk] = PRED35[21];
    PRED35_22_buffer[clk] = PRED35[22];
    PRED35_23_buffer[clk] = PRED35[23];
    PRED35_24_buffer[clk] = PRED35[24];
    PRED35_25_buffer[clk] = PRED35[25];
    PRED35_26_buffer[clk] = PRED35[26];
    PRED35_27_buffer[clk] = PRED35[27];
    PRED35_28_buffer[clk] = PRED35[28];
    PRED35_29_buffer[clk] = PRED35[29];
    PRED35_30_buffer[clk] = PRED35[30];
    PRED35_31_buffer[clk] = PRED35[31];
    PRED36_0_buffer[clk] = PRED36[0];
    PRED36_1_buffer[clk] = PRED36[1];
    PRED36_2_buffer[clk] = PRED36[2];
    PRED36_3_buffer[clk] = PRED36[3];
    PRED36_4_buffer[clk] = PRED36[4];
    PRED36_5_buffer[clk] = PRED36[5];
    PRED36_6_buffer[clk] = PRED36[6];
    PRED36_7_buffer[clk] = PRED36[7];
    PRED36_8_buffer[clk] = PRED36[8];
    PRED36_9_buffer[clk] = PRED36[9];
    PRED36_10_buffer[clk] = PRED36[10];
    PRED36_11_buffer[clk] = PRED36[11];
    PRED36_12_buffer[clk] = PRED36[12];
    PRED36_13_buffer[clk] = PRED36[13];
    PRED36_14_buffer[clk] = PRED36[14];
    PRED36_15_buffer[clk] = PRED36[15];
    PRED36_16_buffer[clk] = PRED36[16];
    PRED36_17_buffer[clk] = PRED36[17];
    PRED36_18_buffer[clk] = PRED36[18];
    PRED36_19_buffer[clk] = PRED36[19];
    PRED36_20_buffer[clk] = PRED36[20];
    PRED36_21_buffer[clk] = PRED36[21];
    PRED36_22_buffer[clk] = PRED36[22];
    PRED36_23_buffer[clk] = PRED36[23];
    PRED36_24_buffer[clk] = PRED36[24];
    PRED36_25_buffer[clk] = PRED36[25];
    PRED36_26_buffer[clk] = PRED36[26];
    PRED36_27_buffer[clk] = PRED36[27];
    PRED36_28_buffer[clk] = PRED36[28];
    PRED36_29_buffer[clk] = PRED36[29];
    PRED36_30_buffer[clk] = PRED36[30];
    PRED36_31_buffer[clk] = PRED36[31];
    PRED37_0_buffer[clk] = PRED37[0];
    PRED37_1_buffer[clk] = PRED37[1];
    PRED37_2_buffer[clk] = PRED37[2];
    PRED37_3_buffer[clk] = PRED37[3];
    PRED37_4_buffer[clk] = PRED37[4];
    PRED37_5_buffer[clk] = PRED37[5];
    PRED37_6_buffer[clk] = PRED37[6];
    PRED37_7_buffer[clk] = PRED37[7];
    PRED37_8_buffer[clk] = PRED37[8];
    PRED37_9_buffer[clk] = PRED37[9];
    PRED37_10_buffer[clk] = PRED37[10];
    PRED37_11_buffer[clk] = PRED37[11];
    PRED37_12_buffer[clk] = PRED37[12];
    PRED37_13_buffer[clk] = PRED37[13];
    PRED37_14_buffer[clk] = PRED37[14];
    PRED37_15_buffer[clk] = PRED37[15];
    PRED37_16_buffer[clk] = PRED37[16];
    PRED37_17_buffer[clk] = PRED37[17];
    PRED37_18_buffer[clk] = PRED37[18];
    PRED37_19_buffer[clk] = PRED37[19];
    PRED37_20_buffer[clk] = PRED37[20];
    PRED37_21_buffer[clk] = PRED37[21];
    PRED37_22_buffer[clk] = PRED37[22];
    PRED37_23_buffer[clk] = PRED37[23];
    PRED37_24_buffer[clk] = PRED37[24];
    PRED37_25_buffer[clk] = PRED37[25];
    PRED37_26_buffer[clk] = PRED37[26];
    PRED37_27_buffer[clk] = PRED37[27];
    PRED37_28_buffer[clk] = PRED37[28];
    PRED37_29_buffer[clk] = PRED37[29];
    PRED37_30_buffer[clk] = PRED37[30];
    PRED37_31_buffer[clk] = PRED37[31];
    PRED38_0_buffer[clk] = PRED38[0];
    PRED38_1_buffer[clk] = PRED38[1];
    PRED38_2_buffer[clk] = PRED38[2];
    PRED38_3_buffer[clk] = PRED38[3];
    PRED38_4_buffer[clk] = PRED38[4];
    PRED38_5_buffer[clk] = PRED38[5];
    PRED38_6_buffer[clk] = PRED38[6];
    PRED38_7_buffer[clk] = PRED38[7];
    PRED38_8_buffer[clk] = PRED38[8];
    PRED38_9_buffer[clk] = PRED38[9];
    PRED38_10_buffer[clk] = PRED38[10];
    PRED38_11_buffer[clk] = PRED38[11];
    PRED38_12_buffer[clk] = PRED38[12];
    PRED38_13_buffer[clk] = PRED38[13];
    PRED38_14_buffer[clk] = PRED38[14];
    PRED38_15_buffer[clk] = PRED38[15];
    PRED38_16_buffer[clk] = PRED38[16];
    PRED38_17_buffer[clk] = PRED38[17];
    PRED38_18_buffer[clk] = PRED38[18];
    PRED38_19_buffer[clk] = PRED38[19];
    PRED38_20_buffer[clk] = PRED38[20];
    PRED38_21_buffer[clk] = PRED38[21];
    PRED38_22_buffer[clk] = PRED38[22];
    PRED38_23_buffer[clk] = PRED38[23];
    PRED38_24_buffer[clk] = PRED38[24];
    PRED38_25_buffer[clk] = PRED38[25];
    PRED38_26_buffer[clk] = PRED38[26];
    PRED38_27_buffer[clk] = PRED38[27];
    PRED38_28_buffer[clk] = PRED38[28];
    PRED38_29_buffer[clk] = PRED38[29];
    PRED38_30_buffer[clk] = PRED38[30];
    PRED38_31_buffer[clk] = PRED38[31];
    PRED39_0_buffer[clk] = PRED39[0];
    PRED39_1_buffer[clk] = PRED39[1];
    PRED39_2_buffer[clk] = PRED39[2];
    PRED39_3_buffer[clk] = PRED39[3];
    PRED39_4_buffer[clk] = PRED39[4];
    PRED39_5_buffer[clk] = PRED39[5];
    PRED39_6_buffer[clk] = PRED39[6];
    PRED39_7_buffer[clk] = PRED39[7];
    PRED39_8_buffer[clk] = PRED39[8];
    PRED39_9_buffer[clk] = PRED39[9];
    PRED39_10_buffer[clk] = PRED39[10];
    PRED39_11_buffer[clk] = PRED39[11];
    PRED39_12_buffer[clk] = PRED39[12];
    PRED39_13_buffer[clk] = PRED39[13];
    PRED39_14_buffer[clk] = PRED39[14];
    PRED39_15_buffer[clk] = PRED39[15];
    PRED39_16_buffer[clk] = PRED39[16];
    PRED39_17_buffer[clk] = PRED39[17];
    PRED39_18_buffer[clk] = PRED39[18];
    PRED39_19_buffer[clk] = PRED39[19];
    PRED39_20_buffer[clk] = PRED39[20];
    PRED39_21_buffer[clk] = PRED39[21];
    PRED39_22_buffer[clk] = PRED39[22];
    PRED39_23_buffer[clk] = PRED39[23];
    PRED39_24_buffer[clk] = PRED39[24];
    PRED39_25_buffer[clk] = PRED39[25];
    PRED39_26_buffer[clk] = PRED39[26];
    PRED39_27_buffer[clk] = PRED39[27];
    PRED39_28_buffer[clk] = PRED39[28];
    PRED39_29_buffer[clk] = PRED39[29];
    PRED39_30_buffer[clk] = PRED39[30];
    PRED39_31_buffer[clk] = PRED39[31];
    PRED40_0_buffer[clk] = PRED40[0];
    PRED40_1_buffer[clk] = PRED40[1];
    PRED40_2_buffer[clk] = PRED40[2];
    PRED40_3_buffer[clk] = PRED40[3];
    PRED40_4_buffer[clk] = PRED40[4];
    PRED40_5_buffer[clk] = PRED40[5];
    PRED40_6_buffer[clk] = PRED40[6];
    PRED40_7_buffer[clk] = PRED40[7];
    PRED40_8_buffer[clk] = PRED40[8];
    PRED40_9_buffer[clk] = PRED40[9];
    PRED40_10_buffer[clk] = PRED40[10];
    PRED40_11_buffer[clk] = PRED40[11];
    PRED40_12_buffer[clk] = PRED40[12];
    PRED40_13_buffer[clk] = PRED40[13];
    PRED40_14_buffer[clk] = PRED40[14];
    PRED40_15_buffer[clk] = PRED40[15];
    PRED40_16_buffer[clk] = PRED40[16];
    PRED40_17_buffer[clk] = PRED40[17];
    PRED40_18_buffer[clk] = PRED40[18];
    PRED40_19_buffer[clk] = PRED40[19];
    PRED40_20_buffer[clk] = PRED40[20];
    PRED40_21_buffer[clk] = PRED40[21];
    PRED40_22_buffer[clk] = PRED40[22];
    PRED40_23_buffer[clk] = PRED40[23];
    PRED40_24_buffer[clk] = PRED40[24];
    PRED40_25_buffer[clk] = PRED40[25];
    PRED40_26_buffer[clk] = PRED40[26];
    PRED40_27_buffer[clk] = PRED40[27];
    PRED40_28_buffer[clk] = PRED40[28];
    PRED40_29_buffer[clk] = PRED40[29];
    PRED40_30_buffer[clk] = PRED40[30];
    PRED40_31_buffer[clk] = PRED40[31];
    PRED41_0_buffer[clk] = PRED41[0];
    PRED41_1_buffer[clk] = PRED41[1];
    PRED41_2_buffer[clk] = PRED41[2];
    PRED41_3_buffer[clk] = PRED41[3];
    PRED41_4_buffer[clk] = PRED41[4];
    PRED41_5_buffer[clk] = PRED41[5];
    PRED41_6_buffer[clk] = PRED41[6];
    PRED41_7_buffer[clk] = PRED41[7];
    PRED41_8_buffer[clk] = PRED41[8];
    PRED41_9_buffer[clk] = PRED41[9];
    PRED41_10_buffer[clk] = PRED41[10];
    PRED41_11_buffer[clk] = PRED41[11];
    PRED41_12_buffer[clk] = PRED41[12];
    PRED41_13_buffer[clk] = PRED41[13];
    PRED41_14_buffer[clk] = PRED41[14];
    PRED41_15_buffer[clk] = PRED41[15];
    PRED41_16_buffer[clk] = PRED41[16];
    PRED41_17_buffer[clk] = PRED41[17];
    PRED41_18_buffer[clk] = PRED41[18];
    PRED41_19_buffer[clk] = PRED41[19];
    PRED41_20_buffer[clk] = PRED41[20];
    PRED41_21_buffer[clk] = PRED41[21];
    PRED41_22_buffer[clk] = PRED41[22];
    PRED41_23_buffer[clk] = PRED41[23];
    PRED41_24_buffer[clk] = PRED41[24];
    PRED41_25_buffer[clk] = PRED41[25];
    PRED41_26_buffer[clk] = PRED41[26];
    PRED41_27_buffer[clk] = PRED41[27];
    PRED41_28_buffer[clk] = PRED41[28];
    PRED41_29_buffer[clk] = PRED41[29];
    PRED41_30_buffer[clk] = PRED41[30];
    PRED41_31_buffer[clk] = PRED41[31];
    PRED42_0_buffer[clk] = PRED42[0];
    PRED42_1_buffer[clk] = PRED42[1];
    PRED42_2_buffer[clk] = PRED42[2];
    PRED42_3_buffer[clk] = PRED42[3];
    PRED42_4_buffer[clk] = PRED42[4];
    PRED42_5_buffer[clk] = PRED42[5];
    PRED42_6_buffer[clk] = PRED42[6];
    PRED42_7_buffer[clk] = PRED42[7];
    PRED42_8_buffer[clk] = PRED42[8];
    PRED42_9_buffer[clk] = PRED42[9];
    PRED42_10_buffer[clk] = PRED42[10];
    PRED42_11_buffer[clk] = PRED42[11];
    PRED42_12_buffer[clk] = PRED42[12];
    PRED42_13_buffer[clk] = PRED42[13];
    PRED42_14_buffer[clk] = PRED42[14];
    PRED42_15_buffer[clk] = PRED42[15];
    PRED42_16_buffer[clk] = PRED42[16];
    PRED42_17_buffer[clk] = PRED42[17];
    PRED42_18_buffer[clk] = PRED42[18];
    PRED42_19_buffer[clk] = PRED42[19];
    PRED42_20_buffer[clk] = PRED42[20];
    PRED42_21_buffer[clk] = PRED42[21];
    PRED42_22_buffer[clk] = PRED42[22];
    PRED42_23_buffer[clk] = PRED42[23];
    PRED42_24_buffer[clk] = PRED42[24];
    PRED42_25_buffer[clk] = PRED42[25];
    PRED42_26_buffer[clk] = PRED42[26];
    PRED42_27_buffer[clk] = PRED42[27];
    PRED42_28_buffer[clk] = PRED42[28];
    PRED42_29_buffer[clk] = PRED42[29];
    PRED42_30_buffer[clk] = PRED42[30];
    PRED42_31_buffer[clk] = PRED42[31];
    PRED43_0_buffer[clk] = PRED43[0];
    PRED43_1_buffer[clk] = PRED43[1];
    PRED43_2_buffer[clk] = PRED43[2];
    PRED43_3_buffer[clk] = PRED43[3];
    PRED43_4_buffer[clk] = PRED43[4];
    PRED43_5_buffer[clk] = PRED43[5];
    PRED43_6_buffer[clk] = PRED43[6];
    PRED43_7_buffer[clk] = PRED43[7];
    PRED43_8_buffer[clk] = PRED43[8];
    PRED43_9_buffer[clk] = PRED43[9];
    PRED43_10_buffer[clk] = PRED43[10];
    PRED43_11_buffer[clk] = PRED43[11];
    PRED43_12_buffer[clk] = PRED43[12];
    PRED43_13_buffer[clk] = PRED43[13];
    PRED43_14_buffer[clk] = PRED43[14];
    PRED43_15_buffer[clk] = PRED43[15];
    PRED43_16_buffer[clk] = PRED43[16];
    PRED43_17_buffer[clk] = PRED43[17];
    PRED43_18_buffer[clk] = PRED43[18];
    PRED43_19_buffer[clk] = PRED43[19];
    PRED43_20_buffer[clk] = PRED43[20];
    PRED43_21_buffer[clk] = PRED43[21];
    PRED43_22_buffer[clk] = PRED43[22];
    PRED43_23_buffer[clk] = PRED43[23];
    PRED43_24_buffer[clk] = PRED43[24];
    PRED43_25_buffer[clk] = PRED43[25];
    PRED43_26_buffer[clk] = PRED43[26];
    PRED43_27_buffer[clk] = PRED43[27];
    PRED43_28_buffer[clk] = PRED43[28];
    PRED43_29_buffer[clk] = PRED43[29];
    PRED43_30_buffer[clk] = PRED43[30];
    PRED43_31_buffer[clk] = PRED43[31];
    PRED44_0_buffer[clk] = PRED44[0];
    PRED44_1_buffer[clk] = PRED44[1];
    PRED44_2_buffer[clk] = PRED44[2];
    PRED44_3_buffer[clk] = PRED44[3];
    PRED44_4_buffer[clk] = PRED44[4];
    PRED44_5_buffer[clk] = PRED44[5];
    PRED44_6_buffer[clk] = PRED44[6];
    PRED44_7_buffer[clk] = PRED44[7];
    PRED44_8_buffer[clk] = PRED44[8];
    PRED44_9_buffer[clk] = PRED44[9];
    PRED44_10_buffer[clk] = PRED44[10];
    PRED44_11_buffer[clk] = PRED44[11];
    PRED44_12_buffer[clk] = PRED44[12];
    PRED44_13_buffer[clk] = PRED44[13];
    PRED44_14_buffer[clk] = PRED44[14];
    PRED44_15_buffer[clk] = PRED44[15];
    PRED44_16_buffer[clk] = PRED44[16];
    PRED44_17_buffer[clk] = PRED44[17];
    PRED44_18_buffer[clk] = PRED44[18];
    PRED44_19_buffer[clk] = PRED44[19];
    PRED44_20_buffer[clk] = PRED44[20];
    PRED44_21_buffer[clk] = PRED44[21];
    PRED44_22_buffer[clk] = PRED44[22];
    PRED44_23_buffer[clk] = PRED44[23];
    PRED44_24_buffer[clk] = PRED44[24];
    PRED44_25_buffer[clk] = PRED44[25];
    PRED44_26_buffer[clk] = PRED44[26];
    PRED44_27_buffer[clk] = PRED44[27];
    PRED44_28_buffer[clk] = PRED44[28];
    PRED44_29_buffer[clk] = PRED44[29];
    PRED44_30_buffer[clk] = PRED44[30];
    PRED44_31_buffer[clk] = PRED44[31];
    PRED45_0_buffer[clk] = PRED45[0];
    PRED45_1_buffer[clk] = PRED45[1];
    PRED45_2_buffer[clk] = PRED45[2];
    PRED45_3_buffer[clk] = PRED45[3];
    PRED45_4_buffer[clk] = PRED45[4];
    PRED45_5_buffer[clk] = PRED45[5];
    PRED45_6_buffer[clk] = PRED45[6];
    PRED45_7_buffer[clk] = PRED45[7];
    PRED45_8_buffer[clk] = PRED45[8];
    PRED45_9_buffer[clk] = PRED45[9];
    PRED45_10_buffer[clk] = PRED45[10];
    PRED45_11_buffer[clk] = PRED45[11];
    PRED45_12_buffer[clk] = PRED45[12];
    PRED45_13_buffer[clk] = PRED45[13];
    PRED45_14_buffer[clk] = PRED45[14];
    PRED45_15_buffer[clk] = PRED45[15];
    PRED45_16_buffer[clk] = PRED45[16];
    PRED45_17_buffer[clk] = PRED45[17];
    PRED45_18_buffer[clk] = PRED45[18];
    PRED45_19_buffer[clk] = PRED45[19];
    PRED45_20_buffer[clk] = PRED45[20];
    PRED45_21_buffer[clk] = PRED45[21];
    PRED45_22_buffer[clk] = PRED45[22];
    PRED45_23_buffer[clk] = PRED45[23];
    PRED45_24_buffer[clk] = PRED45[24];
    PRED45_25_buffer[clk] = PRED45[25];
    PRED45_26_buffer[clk] = PRED45[26];
    PRED45_27_buffer[clk] = PRED45[27];
    PRED45_28_buffer[clk] = PRED45[28];
    PRED45_29_buffer[clk] = PRED45[29];
    PRED45_30_buffer[clk] = PRED45[30];
    PRED45_31_buffer[clk] = PRED45[31];
    PRED46_0_buffer[clk] = PRED46[0];
    PRED46_1_buffer[clk] = PRED46[1];
    PRED46_2_buffer[clk] = PRED46[2];
    PRED46_3_buffer[clk] = PRED46[3];
    PRED46_4_buffer[clk] = PRED46[4];
    PRED46_5_buffer[clk] = PRED46[5];
    PRED46_6_buffer[clk] = PRED46[6];
    PRED46_7_buffer[clk] = PRED46[7];
    PRED46_8_buffer[clk] = PRED46[8];
    PRED46_9_buffer[clk] = PRED46[9];
    PRED46_10_buffer[clk] = PRED46[10];
    PRED46_11_buffer[clk] = PRED46[11];
    PRED46_12_buffer[clk] = PRED46[12];
    PRED46_13_buffer[clk] = PRED46[13];
    PRED46_14_buffer[clk] = PRED46[14];
    PRED46_15_buffer[clk] = PRED46[15];
    PRED46_16_buffer[clk] = PRED46[16];
    PRED46_17_buffer[clk] = PRED46[17];
    PRED46_18_buffer[clk] = PRED46[18];
    PRED46_19_buffer[clk] = PRED46[19];
    PRED46_20_buffer[clk] = PRED46[20];
    PRED46_21_buffer[clk] = PRED46[21];
    PRED46_22_buffer[clk] = PRED46[22];
    PRED46_23_buffer[clk] = PRED46[23];
    PRED46_24_buffer[clk] = PRED46[24];
    PRED46_25_buffer[clk] = PRED46[25];
    PRED46_26_buffer[clk] = PRED46[26];
    PRED46_27_buffer[clk] = PRED46[27];
    PRED46_28_buffer[clk] = PRED46[28];
    PRED46_29_buffer[clk] = PRED46[29];
    PRED46_30_buffer[clk] = PRED46[30];
    PRED46_31_buffer[clk] = PRED46[31];
    PRED47_0_buffer[clk] = PRED47[0];
    PRED47_1_buffer[clk] = PRED47[1];
    PRED47_2_buffer[clk] = PRED47[2];
    PRED47_3_buffer[clk] = PRED47[3];
    PRED47_4_buffer[clk] = PRED47[4];
    PRED47_5_buffer[clk] = PRED47[5];
    PRED47_6_buffer[clk] = PRED47[6];
    PRED47_7_buffer[clk] = PRED47[7];
    PRED47_8_buffer[clk] = PRED47[8];
    PRED47_9_buffer[clk] = PRED47[9];
    PRED47_10_buffer[clk] = PRED47[10];
    PRED47_11_buffer[clk] = PRED47[11];
    PRED47_12_buffer[clk] = PRED47[12];
    PRED47_13_buffer[clk] = PRED47[13];
    PRED47_14_buffer[clk] = PRED47[14];
    PRED47_15_buffer[clk] = PRED47[15];
    PRED47_16_buffer[clk] = PRED47[16];
    PRED47_17_buffer[clk] = PRED47[17];
    PRED47_18_buffer[clk] = PRED47[18];
    PRED47_19_buffer[clk] = PRED47[19];
    PRED47_20_buffer[clk] = PRED47[20];
    PRED47_21_buffer[clk] = PRED47[21];
    PRED47_22_buffer[clk] = PRED47[22];
    PRED47_23_buffer[clk] = PRED47[23];
    PRED47_24_buffer[clk] = PRED47[24];
    PRED47_25_buffer[clk] = PRED47[25];
    PRED47_26_buffer[clk] = PRED47[26];
    PRED47_27_buffer[clk] = PRED47[27];
    PRED47_28_buffer[clk] = PRED47[28];
    PRED47_29_buffer[clk] = PRED47[29];
    PRED47_30_buffer[clk] = PRED47[30];
    PRED47_31_buffer[clk] = PRED47[31];
    PRED48_0_buffer[clk] = PRED48[0];
    PRED48_1_buffer[clk] = PRED48[1];
    PRED48_2_buffer[clk] = PRED48[2];
    PRED48_3_buffer[clk] = PRED48[3];
    PRED48_4_buffer[clk] = PRED48[4];
    PRED48_5_buffer[clk] = PRED48[5];
    PRED48_6_buffer[clk] = PRED48[6];
    PRED48_7_buffer[clk] = PRED48[7];
    PRED48_8_buffer[clk] = PRED48[8];
    PRED48_9_buffer[clk] = PRED48[9];
    PRED48_10_buffer[clk] = PRED48[10];
    PRED48_11_buffer[clk] = PRED48[11];
    PRED48_12_buffer[clk] = PRED48[12];
    PRED48_13_buffer[clk] = PRED48[13];
    PRED48_14_buffer[clk] = PRED48[14];
    PRED48_15_buffer[clk] = PRED48[15];
    PRED48_16_buffer[clk] = PRED48[16];
    PRED48_17_buffer[clk] = PRED48[17];
    PRED48_18_buffer[clk] = PRED48[18];
    PRED48_19_buffer[clk] = PRED48[19];
    PRED48_20_buffer[clk] = PRED48[20];
    PRED48_21_buffer[clk] = PRED48[21];
    PRED48_22_buffer[clk] = PRED48[22];
    PRED48_23_buffer[clk] = PRED48[23];
    PRED48_24_buffer[clk] = PRED48[24];
    PRED48_25_buffer[clk] = PRED48[25];
    PRED48_26_buffer[clk] = PRED48[26];
    PRED48_27_buffer[clk] = PRED48[27];
    PRED48_28_buffer[clk] = PRED48[28];
    PRED48_29_buffer[clk] = PRED48[29];
    PRED48_30_buffer[clk] = PRED48[30];
    PRED48_31_buffer[clk] = PRED48[31];
    PRED49_0_buffer[clk] = PRED49[0];
    PRED49_1_buffer[clk] = PRED49[1];
    PRED49_2_buffer[clk] = PRED49[2];
    PRED49_3_buffer[clk] = PRED49[3];
    PRED49_4_buffer[clk] = PRED49[4];
    PRED49_5_buffer[clk] = PRED49[5];
    PRED49_6_buffer[clk] = PRED49[6];
    PRED49_7_buffer[clk] = PRED49[7];
    PRED49_8_buffer[clk] = PRED49[8];
    PRED49_9_buffer[clk] = PRED49[9];
    PRED49_10_buffer[clk] = PRED49[10];
    PRED49_11_buffer[clk] = PRED49[11];
    PRED49_12_buffer[clk] = PRED49[12];
    PRED49_13_buffer[clk] = PRED49[13];
    PRED49_14_buffer[clk] = PRED49[14];
    PRED49_15_buffer[clk] = PRED49[15];
    PRED49_16_buffer[clk] = PRED49[16];
    PRED49_17_buffer[clk] = PRED49[17];
    PRED49_18_buffer[clk] = PRED49[18];
    PRED49_19_buffer[clk] = PRED49[19];
    PRED49_20_buffer[clk] = PRED49[20];
    PRED49_21_buffer[clk] = PRED49[21];
    PRED49_22_buffer[clk] = PRED49[22];
    PRED49_23_buffer[clk] = PRED49[23];
    PRED49_24_buffer[clk] = PRED49[24];
    PRED49_25_buffer[clk] = PRED49[25];
    PRED49_26_buffer[clk] = PRED49[26];
    PRED49_27_buffer[clk] = PRED49[27];
    PRED49_28_buffer[clk] = PRED49[28];
    PRED49_29_buffer[clk] = PRED49[29];
    PRED49_30_buffer[clk] = PRED49[30];
    PRED49_31_buffer[clk] = PRED49[31];
    PRED50_0_buffer[clk] = PRED50[0];
    PRED50_1_buffer[clk] = PRED50[1];
    PRED50_2_buffer[clk] = PRED50[2];
    PRED50_3_buffer[clk] = PRED50[3];
    PRED50_4_buffer[clk] = PRED50[4];
    PRED50_5_buffer[clk] = PRED50[5];
    PRED50_6_buffer[clk] = PRED50[6];
    PRED50_7_buffer[clk] = PRED50[7];
    PRED50_8_buffer[clk] = PRED50[8];
    PRED50_9_buffer[clk] = PRED50[9];
    PRED50_10_buffer[clk] = PRED50[10];
    PRED50_11_buffer[clk] = PRED50[11];
    PRED50_12_buffer[clk] = PRED50[12];
    PRED50_13_buffer[clk] = PRED50[13];
    PRED50_14_buffer[clk] = PRED50[14];
    PRED50_15_buffer[clk] = PRED50[15];
    PRED50_16_buffer[clk] = PRED50[16];
    PRED50_17_buffer[clk] = PRED50[17];
    PRED50_18_buffer[clk] = PRED50[18];
    PRED50_19_buffer[clk] = PRED50[19];
    PRED50_20_buffer[clk] = PRED50[20];
    PRED50_21_buffer[clk] = PRED50[21];
    PRED50_22_buffer[clk] = PRED50[22];
    PRED50_23_buffer[clk] = PRED50[23];
    PRED50_24_buffer[clk] = PRED50[24];
    PRED50_25_buffer[clk] = PRED50[25];
    PRED50_26_buffer[clk] = PRED50[26];
    PRED50_27_buffer[clk] = PRED50[27];
    PRED50_28_buffer[clk] = PRED50[28];
    PRED50_29_buffer[clk] = PRED50[29];
    PRED50_30_buffer[clk] = PRED50[30];
    PRED50_31_buffer[clk] = PRED50[31];
    PRED51_0_buffer[clk] = PRED51[0];
    PRED51_1_buffer[clk] = PRED51[1];
    PRED51_2_buffer[clk] = PRED51[2];
    PRED51_3_buffer[clk] = PRED51[3];
    PRED51_4_buffer[clk] = PRED51[4];
    PRED51_5_buffer[clk] = PRED51[5];
    PRED51_6_buffer[clk] = PRED51[6];
    PRED51_7_buffer[clk] = PRED51[7];
    PRED51_8_buffer[clk] = PRED51[8];
    PRED51_9_buffer[clk] = PRED51[9];
    PRED51_10_buffer[clk] = PRED51[10];
    PRED51_11_buffer[clk] = PRED51[11];
    PRED51_12_buffer[clk] = PRED51[12];
    PRED51_13_buffer[clk] = PRED51[13];
    PRED51_14_buffer[clk] = PRED51[14];
    PRED51_15_buffer[clk] = PRED51[15];
    PRED51_16_buffer[clk] = PRED51[16];
    PRED51_17_buffer[clk] = PRED51[17];
    PRED51_18_buffer[clk] = PRED51[18];
    PRED51_19_buffer[clk] = PRED51[19];
    PRED51_20_buffer[clk] = PRED51[20];
    PRED51_21_buffer[clk] = PRED51[21];
    PRED51_22_buffer[clk] = PRED51[22];
    PRED51_23_buffer[clk] = PRED51[23];
    PRED51_24_buffer[clk] = PRED51[24];
    PRED51_25_buffer[clk] = PRED51[25];
    PRED51_26_buffer[clk] = PRED51[26];
    PRED51_27_buffer[clk] = PRED51[27];
    PRED51_28_buffer[clk] = PRED51[28];
    PRED51_29_buffer[clk] = PRED51[29];
    PRED51_30_buffer[clk] = PRED51[30];
    PRED51_31_buffer[clk] = PRED51[31];
    PRED52_0_buffer[clk] = PRED52[0];
    PRED52_1_buffer[clk] = PRED52[1];
    PRED52_2_buffer[clk] = PRED52[2];
    PRED52_3_buffer[clk] = PRED52[3];
    PRED52_4_buffer[clk] = PRED52[4];
    PRED52_5_buffer[clk] = PRED52[5];
    PRED52_6_buffer[clk] = PRED52[6];
    PRED52_7_buffer[clk] = PRED52[7];
    PRED52_8_buffer[clk] = PRED52[8];
    PRED52_9_buffer[clk] = PRED52[9];
    PRED52_10_buffer[clk] = PRED52[10];
    PRED52_11_buffer[clk] = PRED52[11];
    PRED52_12_buffer[clk] = PRED52[12];
    PRED52_13_buffer[clk] = PRED52[13];
    PRED52_14_buffer[clk] = PRED52[14];
    PRED52_15_buffer[clk] = PRED52[15];
    PRED52_16_buffer[clk] = PRED52[16];
    PRED52_17_buffer[clk] = PRED52[17];
    PRED52_18_buffer[clk] = PRED52[18];
    PRED52_19_buffer[clk] = PRED52[19];
    PRED52_20_buffer[clk] = PRED52[20];
    PRED52_21_buffer[clk] = PRED52[21];
    PRED52_22_buffer[clk] = PRED52[22];
    PRED52_23_buffer[clk] = PRED52[23];
    PRED52_24_buffer[clk] = PRED52[24];
    PRED52_25_buffer[clk] = PRED52[25];
    PRED52_26_buffer[clk] = PRED52[26];
    PRED52_27_buffer[clk] = PRED52[27];
    PRED52_28_buffer[clk] = PRED52[28];
    PRED52_29_buffer[clk] = PRED52[29];
    PRED52_30_buffer[clk] = PRED52[30];
    PRED52_31_buffer[clk] = PRED52[31];
    PRED53_0_buffer[clk] = PRED53[0];
    PRED53_1_buffer[clk] = PRED53[1];
    PRED53_2_buffer[clk] = PRED53[2];
    PRED53_3_buffer[clk] = PRED53[3];
    PRED53_4_buffer[clk] = PRED53[4];
    PRED53_5_buffer[clk] = PRED53[5];
    PRED53_6_buffer[clk] = PRED53[6];
    PRED53_7_buffer[clk] = PRED53[7];
    PRED53_8_buffer[clk] = PRED53[8];
    PRED53_9_buffer[clk] = PRED53[9];
    PRED53_10_buffer[clk] = PRED53[10];
    PRED53_11_buffer[clk] = PRED53[11];
    PRED53_12_buffer[clk] = PRED53[12];
    PRED53_13_buffer[clk] = PRED53[13];
    PRED53_14_buffer[clk] = PRED53[14];
    PRED53_15_buffer[clk] = PRED53[15];
    PRED53_16_buffer[clk] = PRED53[16];
    PRED53_17_buffer[clk] = PRED53[17];
    PRED53_18_buffer[clk] = PRED53[18];
    PRED53_19_buffer[clk] = PRED53[19];
    PRED53_20_buffer[clk] = PRED53[20];
    PRED53_21_buffer[clk] = PRED53[21];
    PRED53_22_buffer[clk] = PRED53[22];
    PRED53_23_buffer[clk] = PRED53[23];
    PRED53_24_buffer[clk] = PRED53[24];
    PRED53_25_buffer[clk] = PRED53[25];
    PRED53_26_buffer[clk] = PRED53[26];
    PRED53_27_buffer[clk] = PRED53[27];
    PRED53_28_buffer[clk] = PRED53[28];
    PRED53_29_buffer[clk] = PRED53[29];
    PRED53_30_buffer[clk] = PRED53[30];
    PRED53_31_buffer[clk] = PRED53[31];
    PRED54_0_buffer[clk] = PRED54[0];
    PRED54_1_buffer[clk] = PRED54[1];
    PRED54_2_buffer[clk] = PRED54[2];
    PRED54_3_buffer[clk] = PRED54[3];
    PRED54_4_buffer[clk] = PRED54[4];
    PRED54_5_buffer[clk] = PRED54[5];
    PRED54_6_buffer[clk] = PRED54[6];
    PRED54_7_buffer[clk] = PRED54[7];
    PRED54_8_buffer[clk] = PRED54[8];
    PRED54_9_buffer[clk] = PRED54[9];
    PRED54_10_buffer[clk] = PRED54[10];
    PRED54_11_buffer[clk] = PRED54[11];
    PRED54_12_buffer[clk] = PRED54[12];
    PRED54_13_buffer[clk] = PRED54[13];
    PRED54_14_buffer[clk] = PRED54[14];
    PRED54_15_buffer[clk] = PRED54[15];
    PRED54_16_buffer[clk] = PRED54[16];
    PRED54_17_buffer[clk] = PRED54[17];
    PRED54_18_buffer[clk] = PRED54[18];
    PRED54_19_buffer[clk] = PRED54[19];
    PRED54_20_buffer[clk] = PRED54[20];
    PRED54_21_buffer[clk] = PRED54[21];
    PRED54_22_buffer[clk] = PRED54[22];
    PRED54_23_buffer[clk] = PRED54[23];
    PRED54_24_buffer[clk] = PRED54[24];
    PRED54_25_buffer[clk] = PRED54[25];
    PRED54_26_buffer[clk] = PRED54[26];
    PRED54_27_buffer[clk] = PRED54[27];
    PRED54_28_buffer[clk] = PRED54[28];
    PRED54_29_buffer[clk] = PRED54[29];
    PRED54_30_buffer[clk] = PRED54[30];
    PRED54_31_buffer[clk] = PRED54[31];
    PRED55_0_buffer[clk] = PRED55[0];
    PRED55_1_buffer[clk] = PRED55[1];
    PRED55_2_buffer[clk] = PRED55[2];
    PRED55_3_buffer[clk] = PRED55[3];
    PRED55_4_buffer[clk] = PRED55[4];
    PRED55_5_buffer[clk] = PRED55[5];
    PRED55_6_buffer[clk] = PRED55[6];
    PRED55_7_buffer[clk] = PRED55[7];
    PRED55_8_buffer[clk] = PRED55[8];
    PRED55_9_buffer[clk] = PRED55[9];
    PRED55_10_buffer[clk] = PRED55[10];
    PRED55_11_buffer[clk] = PRED55[11];
    PRED55_12_buffer[clk] = PRED55[12];
    PRED55_13_buffer[clk] = PRED55[13];
    PRED55_14_buffer[clk] = PRED55[14];
    PRED55_15_buffer[clk] = PRED55[15];
    PRED55_16_buffer[clk] = PRED55[16];
    PRED55_17_buffer[clk] = PRED55[17];
    PRED55_18_buffer[clk] = PRED55[18];
    PRED55_19_buffer[clk] = PRED55[19];
    PRED55_20_buffer[clk] = PRED55[20];
    PRED55_21_buffer[clk] = PRED55[21];
    PRED55_22_buffer[clk] = PRED55[22];
    PRED55_23_buffer[clk] = PRED55[23];
    PRED55_24_buffer[clk] = PRED55[24];
    PRED55_25_buffer[clk] = PRED55[25];
    PRED55_26_buffer[clk] = PRED55[26];
    PRED55_27_buffer[clk] = PRED55[27];
    PRED55_28_buffer[clk] = PRED55[28];
    PRED55_29_buffer[clk] = PRED55[29];
    PRED55_30_buffer[clk] = PRED55[30];
    PRED55_31_buffer[clk] = PRED55[31];
    PRED56_0_buffer[clk] = PRED56[0];
    PRED56_1_buffer[clk] = PRED56[1];
    PRED56_2_buffer[clk] = PRED56[2];
    PRED56_3_buffer[clk] = PRED56[3];
    PRED56_4_buffer[clk] = PRED56[4];
    PRED56_5_buffer[clk] = PRED56[5];
    PRED56_6_buffer[clk] = PRED56[6];
    PRED56_7_buffer[clk] = PRED56[7];
    PRED56_8_buffer[clk] = PRED56[8];
    PRED56_9_buffer[clk] = PRED56[9];
    PRED56_10_buffer[clk] = PRED56[10];
    PRED56_11_buffer[clk] = PRED56[11];
    PRED56_12_buffer[clk] = PRED56[12];
    PRED56_13_buffer[clk] = PRED56[13];
    PRED56_14_buffer[clk] = PRED56[14];
    PRED56_15_buffer[clk] = PRED56[15];
    PRED56_16_buffer[clk] = PRED56[16];
    PRED56_17_buffer[clk] = PRED56[17];
    PRED56_18_buffer[clk] = PRED56[18];
    PRED56_19_buffer[clk] = PRED56[19];
    PRED56_20_buffer[clk] = PRED56[20];
    PRED56_21_buffer[clk] = PRED56[21];
    PRED56_22_buffer[clk] = PRED56[22];
    PRED56_23_buffer[clk] = PRED56[23];
    PRED56_24_buffer[clk] = PRED56[24];
    PRED56_25_buffer[clk] = PRED56[25];
    PRED56_26_buffer[clk] = PRED56[26];
    PRED56_27_buffer[clk] = PRED56[27];
    PRED56_28_buffer[clk] = PRED56[28];
    PRED56_29_buffer[clk] = PRED56[29];
    PRED56_30_buffer[clk] = PRED56[30];
    PRED56_31_buffer[clk] = PRED56[31];
    PRED57_0_buffer[clk] = PRED57[0];
    PRED57_1_buffer[clk] = PRED57[1];
    PRED57_2_buffer[clk] = PRED57[2];
    PRED57_3_buffer[clk] = PRED57[3];
    PRED57_4_buffer[clk] = PRED57[4];
    PRED57_5_buffer[clk] = PRED57[5];
    PRED57_6_buffer[clk] = PRED57[6];
    PRED57_7_buffer[clk] = PRED57[7];
    PRED57_8_buffer[clk] = PRED57[8];
    PRED57_9_buffer[clk] = PRED57[9];
    PRED57_10_buffer[clk] = PRED57[10];
    PRED57_11_buffer[clk] = PRED57[11];
    PRED57_12_buffer[clk] = PRED57[12];
    PRED57_13_buffer[clk] = PRED57[13];
    PRED57_14_buffer[clk] = PRED57[14];
    PRED57_15_buffer[clk] = PRED57[15];
    PRED57_16_buffer[clk] = PRED57[16];
    PRED57_17_buffer[clk] = PRED57[17];
    PRED57_18_buffer[clk] = PRED57[18];
    PRED57_19_buffer[clk] = PRED57[19];
    PRED57_20_buffer[clk] = PRED57[20];
    PRED57_21_buffer[clk] = PRED57[21];
    PRED57_22_buffer[clk] = PRED57[22];
    PRED57_23_buffer[clk] = PRED57[23];
    PRED57_24_buffer[clk] = PRED57[24];
    PRED57_25_buffer[clk] = PRED57[25];
    PRED57_26_buffer[clk] = PRED57[26];
    PRED57_27_buffer[clk] = PRED57[27];
    PRED57_28_buffer[clk] = PRED57[28];
    PRED57_29_buffer[clk] = PRED57[29];
    PRED57_30_buffer[clk] = PRED57[30];
    PRED57_31_buffer[clk] = PRED57[31];
    PRED58_0_buffer[clk] = PRED58[0];
    PRED58_1_buffer[clk] = PRED58[1];
    PRED58_2_buffer[clk] = PRED58[2];
    PRED58_3_buffer[clk] = PRED58[3];
    PRED58_4_buffer[clk] = PRED58[4];
    PRED58_5_buffer[clk] = PRED58[5];
    PRED58_6_buffer[clk] = PRED58[6];
    PRED58_7_buffer[clk] = PRED58[7];
    PRED58_8_buffer[clk] = PRED58[8];
    PRED58_9_buffer[clk] = PRED58[9];
    PRED58_10_buffer[clk] = PRED58[10];
    PRED58_11_buffer[clk] = PRED58[11];
    PRED58_12_buffer[clk] = PRED58[12];
    PRED58_13_buffer[clk] = PRED58[13];
    PRED58_14_buffer[clk] = PRED58[14];
    PRED58_15_buffer[clk] = PRED58[15];
    PRED58_16_buffer[clk] = PRED58[16];
    PRED58_17_buffer[clk] = PRED58[17];
    PRED58_18_buffer[clk] = PRED58[18];
    PRED58_19_buffer[clk] = PRED58[19];
    PRED58_20_buffer[clk] = PRED58[20];
    PRED58_21_buffer[clk] = PRED58[21];
    PRED58_22_buffer[clk] = PRED58[22];
    PRED58_23_buffer[clk] = PRED58[23];
    PRED58_24_buffer[clk] = PRED58[24];
    PRED58_25_buffer[clk] = PRED58[25];
    PRED58_26_buffer[clk] = PRED58[26];
    PRED58_27_buffer[clk] = PRED58[27];
    PRED58_28_buffer[clk] = PRED58[28];
    PRED58_29_buffer[clk] = PRED58[29];
    PRED58_30_buffer[clk] = PRED58[30];
    PRED58_31_buffer[clk] = PRED58[31];
    PRED59_0_buffer[clk] = PRED59[0];
    PRED59_1_buffer[clk] = PRED59[1];
    PRED59_2_buffer[clk] = PRED59[2];
    PRED59_3_buffer[clk] = PRED59[3];
    PRED59_4_buffer[clk] = PRED59[4];
    PRED59_5_buffer[clk] = PRED59[5];
    PRED59_6_buffer[clk] = PRED59[6];
    PRED59_7_buffer[clk] = PRED59[7];
    PRED59_8_buffer[clk] = PRED59[8];
    PRED59_9_buffer[clk] = PRED59[9];
    PRED59_10_buffer[clk] = PRED59[10];
    PRED59_11_buffer[clk] = PRED59[11];
    PRED59_12_buffer[clk] = PRED59[12];
    PRED59_13_buffer[clk] = PRED59[13];
    PRED59_14_buffer[clk] = PRED59[14];
    PRED59_15_buffer[clk] = PRED59[15];
    PRED59_16_buffer[clk] = PRED59[16];
    PRED59_17_buffer[clk] = PRED59[17];
    PRED59_18_buffer[clk] = PRED59[18];
    PRED59_19_buffer[clk] = PRED59[19];
    PRED59_20_buffer[clk] = PRED59[20];
    PRED59_21_buffer[clk] = PRED59[21];
    PRED59_22_buffer[clk] = PRED59[22];
    PRED59_23_buffer[clk] = PRED59[23];
    PRED59_24_buffer[clk] = PRED59[24];
    PRED59_25_buffer[clk] = PRED59[25];
    PRED59_26_buffer[clk] = PRED59[26];
    PRED59_27_buffer[clk] = PRED59[27];
    PRED59_28_buffer[clk] = PRED59[28];
    PRED59_29_buffer[clk] = PRED59[29];
    PRED59_30_buffer[clk] = PRED59[30];
    PRED59_31_buffer[clk] = PRED59[31];
    PRED60_0_buffer[clk] = PRED60[0];
    PRED60_1_buffer[clk] = PRED60[1];
    PRED60_2_buffer[clk] = PRED60[2];
    PRED60_3_buffer[clk] = PRED60[3];
    PRED60_4_buffer[clk] = PRED60[4];
    PRED60_5_buffer[clk] = PRED60[5];
    PRED60_6_buffer[clk] = PRED60[6];
    PRED60_7_buffer[clk] = PRED60[7];
    PRED60_8_buffer[clk] = PRED60[8];
    PRED60_9_buffer[clk] = PRED60[9];
    PRED60_10_buffer[clk] = PRED60[10];
    PRED60_11_buffer[clk] = PRED60[11];
    PRED60_12_buffer[clk] = PRED60[12];
    PRED60_13_buffer[clk] = PRED60[13];
    PRED60_14_buffer[clk] = PRED60[14];
    PRED60_15_buffer[clk] = PRED60[15];
    PRED60_16_buffer[clk] = PRED60[16];
    PRED60_17_buffer[clk] = PRED60[17];
    PRED60_18_buffer[clk] = PRED60[18];
    PRED60_19_buffer[clk] = PRED60[19];
    PRED60_20_buffer[clk] = PRED60[20];
    PRED60_21_buffer[clk] = PRED60[21];
    PRED60_22_buffer[clk] = PRED60[22];
    PRED60_23_buffer[clk] = PRED60[23];
    PRED60_24_buffer[clk] = PRED60[24];
    PRED60_25_buffer[clk] = PRED60[25];
    PRED60_26_buffer[clk] = PRED60[26];
    PRED60_27_buffer[clk] = PRED60[27];
    PRED60_28_buffer[clk] = PRED60[28];
    PRED60_29_buffer[clk] = PRED60[29];
    PRED60_30_buffer[clk] = PRED60[30];
    PRED60_31_buffer[clk] = PRED60[31];
    PRED61_0_buffer[clk] = PRED61[0];
    PRED61_1_buffer[clk] = PRED61[1];
    PRED61_2_buffer[clk] = PRED61[2];
    PRED61_3_buffer[clk] = PRED61[3];
    PRED61_4_buffer[clk] = PRED61[4];
    PRED61_5_buffer[clk] = PRED61[5];
    PRED61_6_buffer[clk] = PRED61[6];
    PRED61_7_buffer[clk] = PRED61[7];
    PRED61_8_buffer[clk] = PRED61[8];
    PRED61_9_buffer[clk] = PRED61[9];
    PRED61_10_buffer[clk] = PRED61[10];
    PRED61_11_buffer[clk] = PRED61[11];
    PRED61_12_buffer[clk] = PRED61[12];
    PRED61_13_buffer[clk] = PRED61[13];
    PRED61_14_buffer[clk] = PRED61[14];
    PRED61_15_buffer[clk] = PRED61[15];
    PRED61_16_buffer[clk] = PRED61[16];
    PRED61_17_buffer[clk] = PRED61[17];
    PRED61_18_buffer[clk] = PRED61[18];
    PRED61_19_buffer[clk] = PRED61[19];
    PRED61_20_buffer[clk] = PRED61[20];
    PRED61_21_buffer[clk] = PRED61[21];
    PRED61_22_buffer[clk] = PRED61[22];
    PRED61_23_buffer[clk] = PRED61[23];
    PRED61_24_buffer[clk] = PRED61[24];
    PRED61_25_buffer[clk] = PRED61[25];
    PRED61_26_buffer[clk] = PRED61[26];
    PRED61_27_buffer[clk] = PRED61[27];
    PRED61_28_buffer[clk] = PRED61[28];
    PRED61_29_buffer[clk] = PRED61[29];
    PRED61_30_buffer[clk] = PRED61[30];
    PRED61_31_buffer[clk] = PRED61[31];
    PRED62_0_buffer[clk] = PRED62[0];
    PRED62_1_buffer[clk] = PRED62[1];
    PRED62_2_buffer[clk] = PRED62[2];
    PRED62_3_buffer[clk] = PRED62[3];
    PRED62_4_buffer[clk] = PRED62[4];
    PRED62_5_buffer[clk] = PRED62[5];
    PRED62_6_buffer[clk] = PRED62[6];
    PRED62_7_buffer[clk] = PRED62[7];
    PRED62_8_buffer[clk] = PRED62[8];
    PRED62_9_buffer[clk] = PRED62[9];
    PRED62_10_buffer[clk] = PRED62[10];
    PRED62_11_buffer[clk] = PRED62[11];
    PRED62_12_buffer[clk] = PRED62[12];
    PRED62_13_buffer[clk] = PRED62[13];
    PRED62_14_buffer[clk] = PRED62[14];
    PRED62_15_buffer[clk] = PRED62[15];
    PRED62_16_buffer[clk] = PRED62[16];
    PRED62_17_buffer[clk] = PRED62[17];
    PRED62_18_buffer[clk] = PRED62[18];
    PRED62_19_buffer[clk] = PRED62[19];
    PRED62_20_buffer[clk] = PRED62[20];
    PRED62_21_buffer[clk] = PRED62[21];
    PRED62_22_buffer[clk] = PRED62[22];
    PRED62_23_buffer[clk] = PRED62[23];
    PRED62_24_buffer[clk] = PRED62[24];
    PRED62_25_buffer[clk] = PRED62[25];
    PRED62_26_buffer[clk] = PRED62[26];
    PRED62_27_buffer[clk] = PRED62[27];
    PRED62_28_buffer[clk] = PRED62[28];
    PRED62_29_buffer[clk] = PRED62[29];
    PRED62_30_buffer[clk] = PRED62[30];
    PRED62_31_buffer[clk] = PRED62[31];
    PRED63_0_buffer[clk] = PRED63[0];
    PRED63_1_buffer[clk] = PRED63[1];
    PRED63_2_buffer[clk] = PRED63[2];
    PRED63_3_buffer[clk] = PRED63[3];
    PRED63_4_buffer[clk] = PRED63[4];
    PRED63_5_buffer[clk] = PRED63[5];
    PRED63_6_buffer[clk] = PRED63[6];
    PRED63_7_buffer[clk] = PRED63[7];
    PRED63_8_buffer[clk] = PRED63[8];
    PRED63_9_buffer[clk] = PRED63[9];
    PRED63_10_buffer[clk] = PRED63[10];
    PRED63_11_buffer[clk] = PRED63[11];
    PRED63_12_buffer[clk] = PRED63[12];
    PRED63_13_buffer[clk] = PRED63[13];
    PRED63_14_buffer[clk] = PRED63[14];
    PRED63_15_buffer[clk] = PRED63[15];
    PRED63_16_buffer[clk] = PRED63[16];
    PRED63_17_buffer[clk] = PRED63[17];
    PRED63_18_buffer[clk] = PRED63[18];
    PRED63_19_buffer[clk] = PRED63[19];
    PRED63_20_buffer[clk] = PRED63[20];
    PRED63_21_buffer[clk] = PRED63[21];
    PRED63_22_buffer[clk] = PRED63[22];
    PRED63_23_buffer[clk] = PRED63[23];
    PRED63_24_buffer[clk] = PRED63[24];
    PRED63_25_buffer[clk] = PRED63[25];
    PRED63_26_buffer[clk] = PRED63[26];
    PRED63_27_buffer[clk] = PRED63[27];
    PRED63_28_buffer[clk] = PRED63[28];
    PRED63_29_buffer[clk] = PRED63[29];
    PRED63_30_buffer[clk] = PRED63[30];
    PRED63_31_buffer[clk] = PRED63[31];
  end


  // generate warp signal 
  always_comb begin
    if ((PRED0_0_buffer[clk] != PRED0_0_buffer[!clk]) ||(PRED0_1_buffer[clk] != PRED0_1_buffer[!clk]) ||(PRED0_2_buffer[clk] != PRED0_2_buffer[!clk]) ||(PRED0_3_buffer[clk] != PRED0_3_buffer[!clk]) ||(PRED0_4_buffer[clk] != PRED0_4_buffer[!clk]) ||(PRED0_5_buffer[clk] != PRED0_5_buffer[!clk]) ||(PRED0_6_buffer[clk] != PRED0_6_buffer[!clk]) ||(PRED0_7_buffer[clk] != PRED0_7_buffer[!clk]) ||(PRED0_8_buffer[clk] != PRED0_8_buffer[!clk]) ||(PRED0_9_buffer[clk] != PRED0_9_buffer[!clk]) ||(PRED0_10_buffer[clk] != PRED0_10_buffer[!clk]) ||(PRED0_11_buffer[clk] != PRED0_11_buffer[!clk]) ||(PRED0_12_buffer[clk] != PRED0_12_buffer[!clk]) ||(PRED0_13_buffer[clk] != PRED0_13_buffer[!clk]) ||(PRED0_14_buffer[clk] != PRED0_14_buffer[!clk]) ||(PRED0_15_buffer[clk] != PRED0_15_buffer[!clk]) ||(PRED0_16_buffer[clk] != PRED0_16_buffer[!clk]) ||(PRED0_17_buffer[clk] != PRED0_17_buffer[!clk]) ||(PRED0_18_buffer[clk] != PRED0_18_buffer[!clk]) ||(PRED0_19_buffer[clk] != PRED0_19_buffer[!clk]) ||(PRED0_20_buffer[clk] != PRED0_20_buffer[!clk]) ||(PRED0_21_buffer[clk] != PRED0_21_buffer[!clk]) ||(PRED0_22_buffer[clk] != PRED0_22_buffer[!clk]) ||(PRED0_23_buffer[clk] != PRED0_23_buffer[!clk]) ||(PRED0_24_buffer[clk] != PRED0_24_buffer[!clk]) ||(PRED0_25_buffer[clk] != PRED0_25_buffer[!clk]) ||(PRED0_26_buffer[clk] != PRED0_26_buffer[!clk]) ||(PRED0_27_buffer[clk] != PRED0_27_buffer[!clk]) ||(PRED0_28_buffer[clk] != PRED0_28_buffer[!clk]) ||(PRED0_29_buffer[clk] != PRED0_29_buffer[!clk]) ||(PRED0_30_buffer[clk] != PRED0_30_buffer[!clk]) ||(PRED0_31_buffer[clk] != PRED0_31_buffer[!clk]) ||(PRED8_0_buffer[clk] != PRED8_0_buffer[!clk]) ||(PRED8_1_buffer[clk] != PRED8_1_buffer[!clk]) ||(PRED8_2_buffer[clk] != PRED8_2_buffer[!clk]) ||(PRED8_3_buffer[clk] != PRED8_3_buffer[!clk]) ||(PRED8_4_buffer[clk] != PRED8_4_buffer[!clk]) ||(PRED8_5_buffer[clk] != PRED8_5_buffer[!clk]) ||(PRED8_6_buffer[clk] != PRED8_6_buffer[!clk]) ||(PRED8_7_buffer[clk] != PRED8_7_buffer[!clk]) ||(PRED8_8_buffer[clk] != PRED8_8_buffer[!clk]) ||(PRED8_9_buffer[clk] != PRED8_9_buffer[!clk]) ||(PRED8_10_buffer[clk] != PRED8_10_buffer[!clk]) ||(PRED8_11_buffer[clk] != PRED8_11_buffer[!clk]) ||(PRED8_12_buffer[clk] != PRED8_12_buffer[!clk]) ||(PRED8_13_buffer[clk] != PRED8_13_buffer[!clk]) ||(PRED8_14_buffer[clk] != PRED8_14_buffer[!clk]) ||(PRED8_15_buffer[clk] != PRED8_15_buffer[!clk]) ||(PRED8_16_buffer[clk] != PRED8_16_buffer[!clk]) ||(PRED8_17_buffer[clk] != PRED8_17_buffer[!clk]) ||(PRED8_18_buffer[clk] != PRED8_18_buffer[!clk]) ||(PRED8_19_buffer[clk] != PRED8_19_buffer[!clk]) ||(PRED8_20_buffer[clk] != PRED8_20_buffer[!clk]) ||(PRED8_21_buffer[clk] != PRED8_21_buffer[!clk]) ||(PRED8_22_buffer[clk] != PRED8_22_buffer[!clk]) ||(PRED8_23_buffer[clk] != PRED8_23_buffer[!clk]) ||(PRED8_24_buffer[clk] != PRED8_24_buffer[!clk]) ||(PRED8_25_buffer[clk] != PRED8_25_buffer[!clk]) ||(PRED8_26_buffer[clk] != PRED8_26_buffer[!clk]) ||(PRED8_27_buffer[clk] != PRED8_27_buffer[!clk]) ||(PRED8_28_buffer[clk] != PRED8_28_buffer[!clk]) ||(PRED8_29_buffer[clk] != PRED8_29_buffer[!clk]) ||(PRED8_30_buffer[clk] != PRED8_30_buffer[!clk]) ||(PRED8_31_buffer[clk] != PRED8_31_buffer[!clk]) ||(PRED16_0_buffer[clk] != PRED16_0_buffer[!clk]) ||(PRED16_1_buffer[clk] != PRED16_1_buffer[!clk]) ||(PRED16_2_buffer[clk] != PRED16_2_buffer[!clk]) ||(PRED16_3_buffer[clk] != PRED16_3_buffer[!clk]) ||(PRED16_4_buffer[clk] != PRED16_4_buffer[!clk]) ||(PRED16_5_buffer[clk] != PRED16_5_buffer[!clk]) ||(PRED16_6_buffer[clk] != PRED16_6_buffer[!clk]) ||(PRED16_7_buffer[clk] != PRED16_7_buffer[!clk]) ||(PRED16_8_buffer[clk] != PRED16_8_buffer[!clk]) ||(PRED16_9_buffer[clk] != PRED16_9_buffer[!clk]) ||(PRED16_10_buffer[clk] != PRED16_10_buffer[!clk]) ||(PRED16_11_buffer[clk] != PRED16_11_buffer[!clk]) ||(PRED16_12_buffer[clk] != PRED16_12_buffer[!clk]) ||(PRED16_13_buffer[clk] != PRED16_13_buffer[!clk]) ||(PRED16_14_buffer[clk] != PRED16_14_buffer[!clk]) ||(PRED16_15_buffer[clk] != PRED16_15_buffer[!clk]) ||(PRED16_16_buffer[clk] != PRED16_16_buffer[!clk]) ||(PRED16_17_buffer[clk] != PRED16_17_buffer[!clk]) ||(PRED16_18_buffer[clk] != PRED16_18_buffer[!clk]) ||(PRED16_19_buffer[clk] != PRED16_19_buffer[!clk]) ||(PRED16_20_buffer[clk] != PRED16_20_buffer[!clk]) ||(PRED16_21_buffer[clk] != PRED16_21_buffer[!clk]) ||(PRED16_22_buffer[clk] != PRED16_22_buffer[!clk]) ||(PRED16_23_buffer[clk] != PRED16_23_buffer[!clk]) ||(PRED16_24_buffer[clk] != PRED16_24_buffer[!clk]) ||(PRED16_25_buffer[clk] != PRED16_25_buffer[!clk]) ||(PRED16_26_buffer[clk] != PRED16_26_buffer[!clk]) ||(PRED16_27_buffer[clk] != PRED16_27_buffer[!clk]) ||(PRED16_28_buffer[clk] != PRED16_28_buffer[!clk]) ||(PRED16_29_buffer[clk] != PRED16_29_buffer[!clk]) ||(PRED16_30_buffer[clk] != PRED16_30_buffer[!clk]) ||(PRED16_31_buffer[clk] != PRED16_31_buffer[!clk]) ||(PRED24_0_buffer[clk] != PRED24_0_buffer[!clk]) ||(PRED24_1_buffer[clk] != PRED24_1_buffer[!clk]) ||(PRED24_2_buffer[clk] != PRED24_2_buffer[!clk]) ||(PRED24_3_buffer[clk] != PRED24_3_buffer[!clk]) ||(PRED24_4_buffer[clk] != PRED24_4_buffer[!clk]) ||(PRED24_5_buffer[clk] != PRED24_5_buffer[!clk]) ||(PRED24_6_buffer[clk] != PRED24_6_buffer[!clk]) ||(PRED24_7_buffer[clk] != PRED24_7_buffer[!clk]) ||(PRED24_8_buffer[clk] != PRED24_8_buffer[!clk]) ||(PRED24_9_buffer[clk] != PRED24_9_buffer[!clk]) ||(PRED24_10_buffer[clk] != PRED24_10_buffer[!clk]) ||(PRED24_11_buffer[clk] != PRED24_11_buffer[!clk]) ||(PRED24_12_buffer[clk] != PRED24_12_buffer[!clk]) ||(PRED24_13_buffer[clk] != PRED24_13_buffer[!clk]) ||(PRED24_14_buffer[clk] != PRED24_14_buffer[!clk]) ||(PRED24_15_buffer[clk] != PRED24_15_buffer[!clk]) ||(PRED24_16_buffer[clk] != PRED24_16_buffer[!clk]) ||(PRED24_17_buffer[clk] != PRED24_17_buffer[!clk]) ||(PRED24_18_buffer[clk] != PRED24_18_buffer[!clk]) ||(PRED24_19_buffer[clk] != PRED24_19_buffer[!clk]) ||(PRED24_20_buffer[clk] != PRED24_20_buffer[!clk]) ||(PRED24_21_buffer[clk] != PRED24_21_buffer[!clk]) ||(PRED24_22_buffer[clk] != PRED24_22_buffer[!clk]) ||(PRED24_23_buffer[clk] != PRED24_23_buffer[!clk]) ||(PRED24_24_buffer[clk] != PRED24_24_buffer[!clk]) ||(PRED24_25_buffer[clk] != PRED24_25_buffer[!clk]) ||(PRED24_26_buffer[clk] != PRED24_26_buffer[!clk]) ||(PRED24_27_buffer[clk] != PRED24_27_buffer[!clk]) ||(PRED24_28_buffer[clk] != PRED24_28_buffer[!clk]) ||(PRED24_29_buffer[clk] != PRED24_29_buffer[!clk]) ||(PRED24_30_buffer[clk] != PRED24_30_buffer[!clk]) ||(PRED24_31_buffer[clk] != PRED24_31_buffer[!clk]) ||(PRED32_0_buffer[clk] != PRED32_0_buffer[!clk]) ||(PRED32_1_buffer[clk] != PRED32_1_buffer[!clk]) ||(PRED32_2_buffer[clk] != PRED32_2_buffer[!clk]) ||(PRED32_3_buffer[clk] != PRED32_3_buffer[!clk]) ||(PRED32_4_buffer[clk] != PRED32_4_buffer[!clk]) ||(PRED32_5_buffer[clk] != PRED32_5_buffer[!clk]) ||(PRED32_6_buffer[clk] != PRED32_6_buffer[!clk]) ||(PRED32_7_buffer[clk] != PRED32_7_buffer[!clk]) ||(PRED32_8_buffer[clk] != PRED32_8_buffer[!clk]) ||(PRED32_9_buffer[clk] != PRED32_9_buffer[!clk]) ||(PRED32_10_buffer[clk] != PRED32_10_buffer[!clk]) ||(PRED32_11_buffer[clk] != PRED32_11_buffer[!clk]) ||(PRED32_12_buffer[clk] != PRED32_12_buffer[!clk]) ||(PRED32_13_buffer[clk] != PRED32_13_buffer[!clk]) ||(PRED32_14_buffer[clk] != PRED32_14_buffer[!clk]) ||(PRED32_15_buffer[clk] != PRED32_15_buffer[!clk]) ||(PRED32_16_buffer[clk] != PRED32_16_buffer[!clk]) ||(PRED32_17_buffer[clk] != PRED32_17_buffer[!clk]) ||(PRED32_18_buffer[clk] != PRED32_18_buffer[!clk]) ||(PRED32_19_buffer[clk] != PRED32_19_buffer[!clk]) ||(PRED32_20_buffer[clk] != PRED32_20_buffer[!clk]) ||(PRED32_21_buffer[clk] != PRED32_21_buffer[!clk]) ||(PRED32_22_buffer[clk] != PRED32_22_buffer[!clk]) ||(PRED32_23_buffer[clk] != PRED32_23_buffer[!clk]) ||(PRED32_24_buffer[clk] != PRED32_24_buffer[!clk]) ||(PRED32_25_buffer[clk] != PRED32_25_buffer[!clk]) ||(PRED32_26_buffer[clk] != PRED32_26_buffer[!clk]) ||(PRED32_27_buffer[clk] != PRED32_27_buffer[!clk]) ||(PRED32_28_buffer[clk] != PRED32_28_buffer[!clk]) ||(PRED32_29_buffer[clk] != PRED32_29_buffer[!clk]) ||(PRED32_30_buffer[clk] != PRED32_30_buffer[!clk]) ||(PRED32_31_buffer[clk] != PRED32_31_buffer[!clk]) ||(PRED40_0_buffer[clk] != PRED40_0_buffer[!clk]) ||(PRED40_1_buffer[clk] != PRED40_1_buffer[!clk]) ||(PRED40_2_buffer[clk] != PRED40_2_buffer[!clk]) ||(PRED40_3_buffer[clk] != PRED40_3_buffer[!clk]) ||(PRED40_4_buffer[clk] != PRED40_4_buffer[!clk]) ||(PRED40_5_buffer[clk] != PRED40_5_buffer[!clk]) ||(PRED40_6_buffer[clk] != PRED40_6_buffer[!clk]) ||(PRED40_7_buffer[clk] != PRED40_7_buffer[!clk]) ||(PRED40_8_buffer[clk] != PRED40_8_buffer[!clk]) ||(PRED40_9_buffer[clk] != PRED40_9_buffer[!clk]) ||(PRED40_10_buffer[clk] != PRED40_10_buffer[!clk]) ||(PRED40_11_buffer[clk] != PRED40_11_buffer[!clk]) ||(PRED40_12_buffer[clk] != PRED40_12_buffer[!clk]) ||(PRED40_13_buffer[clk] != PRED40_13_buffer[!clk]) ||(PRED40_14_buffer[clk] != PRED40_14_buffer[!clk]) ||(PRED40_15_buffer[clk] != PRED40_15_buffer[!clk]) ||(PRED40_16_buffer[clk] != PRED40_16_buffer[!clk]) ||(PRED40_17_buffer[clk] != PRED40_17_buffer[!clk]) ||(PRED40_18_buffer[clk] != PRED40_18_buffer[!clk]) ||(PRED40_19_buffer[clk] != PRED40_19_buffer[!clk]) ||(PRED40_20_buffer[clk] != PRED40_20_buffer[!clk]) ||(PRED40_21_buffer[clk] != PRED40_21_buffer[!clk]) ||(PRED40_22_buffer[clk] != PRED40_22_buffer[!clk]) ||(PRED40_23_buffer[clk] != PRED40_23_buffer[!clk]) ||(PRED40_24_buffer[clk] != PRED40_24_buffer[!clk]) ||(PRED40_25_buffer[clk] != PRED40_25_buffer[!clk]) ||(PRED40_26_buffer[clk] != PRED40_26_buffer[!clk]) ||(PRED40_27_buffer[clk] != PRED40_27_buffer[!clk]) ||(PRED40_28_buffer[clk] != PRED40_28_buffer[!clk]) ||(PRED40_29_buffer[clk] != PRED40_29_buffer[!clk]) ||(PRED40_30_buffer[clk] != PRED40_30_buffer[!clk]) ||(PRED40_31_buffer[clk] != PRED40_31_buffer[!clk]) ||(PRED48_0_buffer[clk] != PRED48_0_buffer[!clk]) ||(PRED48_1_buffer[clk] != PRED48_1_buffer[!clk]) ||(PRED48_2_buffer[clk] != PRED48_2_buffer[!clk]) ||(PRED48_3_buffer[clk] != PRED48_3_buffer[!clk]) ||(PRED48_4_buffer[clk] != PRED48_4_buffer[!clk]) ||(PRED48_5_buffer[clk] != PRED48_5_buffer[!clk]) ||(PRED48_6_buffer[clk] != PRED48_6_buffer[!clk]) ||(PRED48_7_buffer[clk] != PRED48_7_buffer[!clk]) ||(PRED48_8_buffer[clk] != PRED48_8_buffer[!clk]) ||(PRED48_9_buffer[clk] != PRED48_9_buffer[!clk]) ||(PRED48_10_buffer[clk] != PRED48_10_buffer[!clk]) ||(PRED48_11_buffer[clk] != PRED48_11_buffer[!clk]) ||(PRED48_12_buffer[clk] != PRED48_12_buffer[!clk]) ||(PRED48_13_buffer[clk] != PRED48_13_buffer[!clk]) ||(PRED48_14_buffer[clk] != PRED48_14_buffer[!clk]) ||(PRED48_15_buffer[clk] != PRED48_15_buffer[!clk]) ||(PRED48_16_buffer[clk] != PRED48_16_buffer[!clk]) ||(PRED48_17_buffer[clk] != PRED48_17_buffer[!clk]) ||(PRED48_18_buffer[clk] != PRED48_18_buffer[!clk]) ||(PRED48_19_buffer[clk] != PRED48_19_buffer[!clk]) ||(PRED48_20_buffer[clk] != PRED48_20_buffer[!clk]) ||(PRED48_21_buffer[clk] != PRED48_21_buffer[!clk]) ||(PRED48_22_buffer[clk] != PRED48_22_buffer[!clk]) ||(PRED48_23_buffer[clk] != PRED48_23_buffer[!clk]) ||(PRED48_24_buffer[clk] != PRED48_24_buffer[!clk]) ||(PRED48_25_buffer[clk] != PRED48_25_buffer[!clk]) ||(PRED48_26_buffer[clk] != PRED48_26_buffer[!clk]) ||(PRED48_27_buffer[clk] != PRED48_27_buffer[!clk]) ||(PRED48_28_buffer[clk] != PRED48_28_buffer[!clk]) ||(PRED48_29_buffer[clk] != PRED48_29_buffer[!clk]) ||(PRED48_30_buffer[clk] != PRED48_30_buffer[!clk]) ||(PRED48_31_buffer[clk] != PRED48_31_buffer[!clk]) ||(PRED56_0_buffer[clk] != PRED56_0_buffer[!clk]) ||(PRED56_1_buffer[clk] != PRED56_1_buffer[!clk]) ||(PRED56_2_buffer[clk] != PRED56_2_buffer[!clk]) ||(PRED56_3_buffer[clk] != PRED56_3_buffer[!clk]) ||(PRED56_4_buffer[clk] != PRED56_4_buffer[!clk]) ||(PRED56_5_buffer[clk] != PRED56_5_buffer[!clk]) ||(PRED56_6_buffer[clk] != PRED56_6_buffer[!clk]) ||(PRED56_7_buffer[clk] != PRED56_7_buffer[!clk]) ||(PRED56_8_buffer[clk] != PRED56_8_buffer[!clk]) ||(PRED56_9_buffer[clk] != PRED56_9_buffer[!clk]) ||(PRED56_10_buffer[clk] != PRED56_10_buffer[!clk]) ||(PRED56_11_buffer[clk] != PRED56_11_buffer[!clk]) ||(PRED56_12_buffer[clk] != PRED56_12_buffer[!clk]) ||(PRED56_13_buffer[clk] != PRED56_13_buffer[!clk]) ||(PRED56_14_buffer[clk] != PRED56_14_buffer[!clk]) ||(PRED56_15_buffer[clk] != PRED56_15_buffer[!clk]) ||(PRED56_16_buffer[clk] != PRED56_16_buffer[!clk]) ||(PRED56_17_buffer[clk] != PRED56_17_buffer[!clk]) ||(PRED56_18_buffer[clk] != PRED56_18_buffer[!clk]) ||(PRED56_19_buffer[clk] != PRED56_19_buffer[!clk]) ||(PRED56_20_buffer[clk] != PRED56_20_buffer[!clk]) ||(PRED56_21_buffer[clk] != PRED56_21_buffer[!clk]) ||(PRED56_22_buffer[clk] != PRED56_22_buffer[!clk]) ||(PRED56_23_buffer[clk] != PRED56_23_buffer[!clk]) ||(PRED56_24_buffer[clk] != PRED56_24_buffer[!clk]) ||(PRED56_25_buffer[clk] != PRED56_25_buffer[!clk]) ||(PRED56_26_buffer[clk] != PRED56_26_buffer[!clk]) ||(PRED56_27_buffer[clk] != PRED56_27_buffer[!clk]) ||(PRED56_28_buffer[clk] != PRED56_28_buffer[!clk]) ||(PRED56_29_buffer[clk] != PRED56_29_buffer[!clk]) ||(PRED56_30_buffer[clk] != PRED56_30_buffer[!clk]) ||(PRED56_31_buffer[clk] != PRED56_31_buffer[!clk]) ) begin
      warp0_sig = 1'b1;
    end else begin
      warp0_sig = 1'b0;
    end

    if ((PRED1_0_buffer[clk] != PRED1_0_buffer[!clk]) ||(PRED1_1_buffer[clk] != PRED1_1_buffer[!clk]) ||(PRED1_2_buffer[clk] != PRED1_2_buffer[!clk]) ||(PRED1_3_buffer[clk] != PRED1_3_buffer[!clk]) ||(PRED1_4_buffer[clk] != PRED1_4_buffer[!clk]) ||(PRED1_5_buffer[clk] != PRED1_5_buffer[!clk]) ||(PRED1_6_buffer[clk] != PRED1_6_buffer[!clk]) ||(PRED1_7_buffer[clk] != PRED1_7_buffer[!clk]) ||(PRED1_8_buffer[clk] != PRED1_8_buffer[!clk]) ||(PRED1_9_buffer[clk] != PRED1_9_buffer[!clk]) ||(PRED1_10_buffer[clk] != PRED1_10_buffer[!clk]) ||(PRED1_11_buffer[clk] != PRED1_11_buffer[!clk]) ||(PRED1_12_buffer[clk] != PRED1_12_buffer[!clk]) ||(PRED1_13_buffer[clk] != PRED1_13_buffer[!clk]) ||(PRED1_14_buffer[clk] != PRED1_14_buffer[!clk]) ||(PRED1_15_buffer[clk] != PRED1_15_buffer[!clk]) ||(PRED1_16_buffer[clk] != PRED1_16_buffer[!clk]) ||(PRED1_17_buffer[clk] != PRED1_17_buffer[!clk]) ||(PRED1_18_buffer[clk] != PRED1_18_buffer[!clk]) ||(PRED1_19_buffer[clk] != PRED1_19_buffer[!clk]) ||(PRED1_20_buffer[clk] != PRED1_20_buffer[!clk]) ||(PRED1_21_buffer[clk] != PRED1_21_buffer[!clk]) ||(PRED1_22_buffer[clk] != PRED1_22_buffer[!clk]) ||(PRED1_23_buffer[clk] != PRED1_23_buffer[!clk]) ||(PRED1_24_buffer[clk] != PRED1_24_buffer[!clk]) ||(PRED1_25_buffer[clk] != PRED1_25_buffer[!clk]) ||(PRED1_26_buffer[clk] != PRED1_26_buffer[!clk]) ||(PRED1_27_buffer[clk] != PRED1_27_buffer[!clk]) ||(PRED1_28_buffer[clk] != PRED1_28_buffer[!clk]) ||(PRED1_29_buffer[clk] != PRED1_29_buffer[!clk]) ||(PRED1_30_buffer[clk] != PRED1_30_buffer[!clk]) ||(PRED1_31_buffer[clk] != PRED1_31_buffer[!clk]) ||(PRED9_0_buffer[clk] != PRED9_0_buffer[!clk]) ||(PRED9_1_buffer[clk] != PRED9_1_buffer[!clk]) ||(PRED9_2_buffer[clk] != PRED9_2_buffer[!clk]) ||(PRED9_3_buffer[clk] != PRED9_3_buffer[!clk]) ||(PRED9_4_buffer[clk] != PRED9_4_buffer[!clk]) ||(PRED9_5_buffer[clk] != PRED9_5_buffer[!clk]) ||(PRED9_6_buffer[clk] != PRED9_6_buffer[!clk]) ||(PRED9_7_buffer[clk] != PRED9_7_buffer[!clk]) ||(PRED9_8_buffer[clk] != PRED9_8_buffer[!clk]) ||(PRED9_9_buffer[clk] != PRED9_9_buffer[!clk]) ||(PRED9_10_buffer[clk] != PRED9_10_buffer[!clk]) ||(PRED9_11_buffer[clk] != PRED9_11_buffer[!clk]) ||(PRED9_12_buffer[clk] != PRED9_12_buffer[!clk]) ||(PRED9_13_buffer[clk] != PRED9_13_buffer[!clk]) ||(PRED9_14_buffer[clk] != PRED9_14_buffer[!clk]) ||(PRED9_15_buffer[clk] != PRED9_15_buffer[!clk]) ||(PRED9_16_buffer[clk] != PRED9_16_buffer[!clk]) ||(PRED9_17_buffer[clk] != PRED9_17_buffer[!clk]) ||(PRED9_18_buffer[clk] != PRED9_18_buffer[!clk]) ||(PRED9_19_buffer[clk] != PRED9_19_buffer[!clk]) ||(PRED9_20_buffer[clk] != PRED9_20_buffer[!clk]) ||(PRED9_21_buffer[clk] != PRED9_21_buffer[!clk]) ||(PRED9_22_buffer[clk] != PRED9_22_buffer[!clk]) ||(PRED9_23_buffer[clk] != PRED9_23_buffer[!clk]) ||(PRED9_24_buffer[clk] != PRED9_24_buffer[!clk]) ||(PRED9_25_buffer[clk] != PRED9_25_buffer[!clk]) ||(PRED9_26_buffer[clk] != PRED9_26_buffer[!clk]) ||(PRED9_27_buffer[clk] != PRED9_27_buffer[!clk]) ||(PRED9_28_buffer[clk] != PRED9_28_buffer[!clk]) ||(PRED9_29_buffer[clk] != PRED9_29_buffer[!clk]) ||(PRED9_30_buffer[clk] != PRED9_30_buffer[!clk]) ||(PRED9_31_buffer[clk] != PRED9_31_buffer[!clk]) ||(PRED17_0_buffer[clk] != PRED17_0_buffer[!clk]) ||(PRED17_1_buffer[clk] != PRED17_1_buffer[!clk]) ||(PRED17_2_buffer[clk] != PRED17_2_buffer[!clk]) ||(PRED17_3_buffer[clk] != PRED17_3_buffer[!clk]) ||(PRED17_4_buffer[clk] != PRED17_4_buffer[!clk]) ||(PRED17_5_buffer[clk] != PRED17_5_buffer[!clk]) ||(PRED17_6_buffer[clk] != PRED17_6_buffer[!clk]) ||(PRED17_7_buffer[clk] != PRED17_7_buffer[!clk]) ||(PRED17_8_buffer[clk] != PRED17_8_buffer[!clk]) ||(PRED17_9_buffer[clk] != PRED17_9_buffer[!clk]) ||(PRED17_10_buffer[clk] != PRED17_10_buffer[!clk]) ||(PRED17_11_buffer[clk] != PRED17_11_buffer[!clk]) ||(PRED17_12_buffer[clk] != PRED17_12_buffer[!clk]) ||(PRED17_13_buffer[clk] != PRED17_13_buffer[!clk]) ||(PRED17_14_buffer[clk] != PRED17_14_buffer[!clk]) ||(PRED17_15_buffer[clk] != PRED17_15_buffer[!clk]) ||(PRED17_16_buffer[clk] != PRED17_16_buffer[!clk]) ||(PRED17_17_buffer[clk] != PRED17_17_buffer[!clk]) ||(PRED17_18_buffer[clk] != PRED17_18_buffer[!clk]) ||(PRED17_19_buffer[clk] != PRED17_19_buffer[!clk]) ||(PRED17_20_buffer[clk] != PRED17_20_buffer[!clk]) ||(PRED17_21_buffer[clk] != PRED17_21_buffer[!clk]) ||(PRED17_22_buffer[clk] != PRED17_22_buffer[!clk]) ||(PRED17_23_buffer[clk] != PRED17_23_buffer[!clk]) ||(PRED17_24_buffer[clk] != PRED17_24_buffer[!clk]) ||(PRED17_25_buffer[clk] != PRED17_25_buffer[!clk]) ||(PRED17_26_buffer[clk] != PRED17_26_buffer[!clk]) ||(PRED17_27_buffer[clk] != PRED17_27_buffer[!clk]) ||(PRED17_28_buffer[clk] != PRED17_28_buffer[!clk]) ||(PRED17_29_buffer[clk] != PRED17_29_buffer[!clk]) ||(PRED17_30_buffer[clk] != PRED17_30_buffer[!clk]) ||(PRED17_31_buffer[clk] != PRED17_31_buffer[!clk]) ||(PRED25_0_buffer[clk] != PRED25_0_buffer[!clk]) ||(PRED25_1_buffer[clk] != PRED25_1_buffer[!clk]) ||(PRED25_2_buffer[clk] != PRED25_2_buffer[!clk]) ||(PRED25_3_buffer[clk] != PRED25_3_buffer[!clk]) ||(PRED25_4_buffer[clk] != PRED25_4_buffer[!clk]) ||(PRED25_5_buffer[clk] != PRED25_5_buffer[!clk]) ||(PRED25_6_buffer[clk] != PRED25_6_buffer[!clk]) ||(PRED25_7_buffer[clk] != PRED25_7_buffer[!clk]) ||(PRED25_8_buffer[clk] != PRED25_8_buffer[!clk]) ||(PRED25_9_buffer[clk] != PRED25_9_buffer[!clk]) ||(PRED25_10_buffer[clk] != PRED25_10_buffer[!clk]) ||(PRED25_11_buffer[clk] != PRED25_11_buffer[!clk]) ||(PRED25_12_buffer[clk] != PRED25_12_buffer[!clk]) ||(PRED25_13_buffer[clk] != PRED25_13_buffer[!clk]) ||(PRED25_14_buffer[clk] != PRED25_14_buffer[!clk]) ||(PRED25_15_buffer[clk] != PRED25_15_buffer[!clk]) ||(PRED25_16_buffer[clk] != PRED25_16_buffer[!clk]) ||(PRED25_17_buffer[clk] != PRED25_17_buffer[!clk]) ||(PRED25_18_buffer[clk] != PRED25_18_buffer[!clk]) ||(PRED25_19_buffer[clk] != PRED25_19_buffer[!clk]) ||(PRED25_20_buffer[clk] != PRED25_20_buffer[!clk]) ||(PRED25_21_buffer[clk] != PRED25_21_buffer[!clk]) ||(PRED25_22_buffer[clk] != PRED25_22_buffer[!clk]) ||(PRED25_23_buffer[clk] != PRED25_23_buffer[!clk]) ||(PRED25_24_buffer[clk] != PRED25_24_buffer[!clk]) ||(PRED25_25_buffer[clk] != PRED25_25_buffer[!clk]) ||(PRED25_26_buffer[clk] != PRED25_26_buffer[!clk]) ||(PRED25_27_buffer[clk] != PRED25_27_buffer[!clk]) ||(PRED25_28_buffer[clk] != PRED25_28_buffer[!clk]) ||(PRED25_29_buffer[clk] != PRED25_29_buffer[!clk]) ||(PRED25_30_buffer[clk] != PRED25_30_buffer[!clk]) ||(PRED25_31_buffer[clk] != PRED25_31_buffer[!clk]) ||(PRED33_0_buffer[clk] != PRED33_0_buffer[!clk]) ||(PRED33_1_buffer[clk] != PRED33_1_buffer[!clk]) ||(PRED33_2_buffer[clk] != PRED33_2_buffer[!clk]) ||(PRED33_3_buffer[clk] != PRED33_3_buffer[!clk]) ||(PRED33_4_buffer[clk] != PRED33_4_buffer[!clk]) ||(PRED33_5_buffer[clk] != PRED33_5_buffer[!clk]) ||(PRED33_6_buffer[clk] != PRED33_6_buffer[!clk]) ||(PRED33_7_buffer[clk] != PRED33_7_buffer[!clk]) ||(PRED33_8_buffer[clk] != PRED33_8_buffer[!clk]) ||(PRED33_9_buffer[clk] != PRED33_9_buffer[!clk]) ||(PRED33_10_buffer[clk] != PRED33_10_buffer[!clk]) ||(PRED33_11_buffer[clk] != PRED33_11_buffer[!clk]) ||(PRED33_12_buffer[clk] != PRED33_12_buffer[!clk]) ||(PRED33_13_buffer[clk] != PRED33_13_buffer[!clk]) ||(PRED33_14_buffer[clk] != PRED33_14_buffer[!clk]) ||(PRED33_15_buffer[clk] != PRED33_15_buffer[!clk]) ||(PRED33_16_buffer[clk] != PRED33_16_buffer[!clk]) ||(PRED33_17_buffer[clk] != PRED33_17_buffer[!clk]) ||(PRED33_18_buffer[clk] != PRED33_18_buffer[!clk]) ||(PRED33_19_buffer[clk] != PRED33_19_buffer[!clk]) ||(PRED33_20_buffer[clk] != PRED33_20_buffer[!clk]) ||(PRED33_21_buffer[clk] != PRED33_21_buffer[!clk]) ||(PRED33_22_buffer[clk] != PRED33_22_buffer[!clk]) ||(PRED33_23_buffer[clk] != PRED33_23_buffer[!clk]) ||(PRED33_24_buffer[clk] != PRED33_24_buffer[!clk]) ||(PRED33_25_buffer[clk] != PRED33_25_buffer[!clk]) ||(PRED33_26_buffer[clk] != PRED33_26_buffer[!clk]) ||(PRED33_27_buffer[clk] != PRED33_27_buffer[!clk]) ||(PRED33_28_buffer[clk] != PRED33_28_buffer[!clk]) ||(PRED33_29_buffer[clk] != PRED33_29_buffer[!clk]) ||(PRED33_30_buffer[clk] != PRED33_30_buffer[!clk]) ||(PRED33_31_buffer[clk] != PRED33_31_buffer[!clk]) ||(PRED41_0_buffer[clk] != PRED41_0_buffer[!clk]) ||(PRED41_1_buffer[clk] != PRED41_1_buffer[!clk]) ||(PRED41_2_buffer[clk] != PRED41_2_buffer[!clk]) ||(PRED41_3_buffer[clk] != PRED41_3_buffer[!clk]) ||(PRED41_4_buffer[clk] != PRED41_4_buffer[!clk]) ||(PRED41_5_buffer[clk] != PRED41_5_buffer[!clk]) ||(PRED41_6_buffer[clk] != PRED41_6_buffer[!clk]) ||(PRED41_7_buffer[clk] != PRED41_7_buffer[!clk]) ||(PRED41_8_buffer[clk] != PRED41_8_buffer[!clk]) ||(PRED41_9_buffer[clk] != PRED41_9_buffer[!clk]) ||(PRED41_10_buffer[clk] != PRED41_10_buffer[!clk]) ||(PRED41_11_buffer[clk] != PRED41_11_buffer[!clk]) ||(PRED41_12_buffer[clk] != PRED41_12_buffer[!clk]) ||(PRED41_13_buffer[clk] != PRED41_13_buffer[!clk]) ||(PRED41_14_buffer[clk] != PRED41_14_buffer[!clk]) ||(PRED41_15_buffer[clk] != PRED41_15_buffer[!clk]) ||(PRED41_16_buffer[clk] != PRED41_16_buffer[!clk]) ||(PRED41_17_buffer[clk] != PRED41_17_buffer[!clk]) ||(PRED41_18_buffer[clk] != PRED41_18_buffer[!clk]) ||(PRED41_19_buffer[clk] != PRED41_19_buffer[!clk]) ||(PRED41_20_buffer[clk] != PRED41_20_buffer[!clk]) ||(PRED41_21_buffer[clk] != PRED41_21_buffer[!clk]) ||(PRED41_22_buffer[clk] != PRED41_22_buffer[!clk]) ||(PRED41_23_buffer[clk] != PRED41_23_buffer[!clk]) ||(PRED41_24_buffer[clk] != PRED41_24_buffer[!clk]) ||(PRED41_25_buffer[clk] != PRED41_25_buffer[!clk]) ||(PRED41_26_buffer[clk] != PRED41_26_buffer[!clk]) ||(PRED41_27_buffer[clk] != PRED41_27_buffer[!clk]) ||(PRED41_28_buffer[clk] != PRED41_28_buffer[!clk]) ||(PRED41_29_buffer[clk] != PRED41_29_buffer[!clk]) ||(PRED41_30_buffer[clk] != PRED41_30_buffer[!clk]) ||(PRED41_31_buffer[clk] != PRED41_31_buffer[!clk]) ||(PRED49_0_buffer[clk] != PRED49_0_buffer[!clk]) ||(PRED49_1_buffer[clk] != PRED49_1_buffer[!clk]) ||(PRED49_2_buffer[clk] != PRED49_2_buffer[!clk]) ||(PRED49_3_buffer[clk] != PRED49_3_buffer[!clk]) ||(PRED49_4_buffer[clk] != PRED49_4_buffer[!clk]) ||(PRED49_5_buffer[clk] != PRED49_5_buffer[!clk]) ||(PRED49_6_buffer[clk] != PRED49_6_buffer[!clk]) ||(PRED49_7_buffer[clk] != PRED49_7_buffer[!clk]) ||(PRED49_8_buffer[clk] != PRED49_8_buffer[!clk]) ||(PRED49_9_buffer[clk] != PRED49_9_buffer[!clk]) ||(PRED49_10_buffer[clk] != PRED49_10_buffer[!clk]) ||(PRED49_11_buffer[clk] != PRED49_11_buffer[!clk]) ||(PRED49_12_buffer[clk] != PRED49_12_buffer[!clk]) ||(PRED49_13_buffer[clk] != PRED49_13_buffer[!clk]) ||(PRED49_14_buffer[clk] != PRED49_14_buffer[!clk]) ||(PRED49_15_buffer[clk] != PRED49_15_buffer[!clk]) ||(PRED49_16_buffer[clk] != PRED49_16_buffer[!clk]) ||(PRED49_17_buffer[clk] != PRED49_17_buffer[!clk]) ||(PRED49_18_buffer[clk] != PRED49_18_buffer[!clk]) ||(PRED49_19_buffer[clk] != PRED49_19_buffer[!clk]) ||(PRED49_20_buffer[clk] != PRED49_20_buffer[!clk]) ||(PRED49_21_buffer[clk] != PRED49_21_buffer[!clk]) ||(PRED49_22_buffer[clk] != PRED49_22_buffer[!clk]) ||(PRED49_23_buffer[clk] != PRED49_23_buffer[!clk]) ||(PRED49_24_buffer[clk] != PRED49_24_buffer[!clk]) ||(PRED49_25_buffer[clk] != PRED49_25_buffer[!clk]) ||(PRED49_26_buffer[clk] != PRED49_26_buffer[!clk]) ||(PRED49_27_buffer[clk] != PRED49_27_buffer[!clk]) ||(PRED49_28_buffer[clk] != PRED49_28_buffer[!clk]) ||(PRED49_29_buffer[clk] != PRED49_29_buffer[!clk]) ||(PRED49_30_buffer[clk] != PRED49_30_buffer[!clk]) ||(PRED49_31_buffer[clk] != PRED49_31_buffer[!clk]) ||(PRED57_0_buffer[clk] != PRED57_0_buffer[!clk]) ||(PRED57_1_buffer[clk] != PRED57_1_buffer[!clk]) ||(PRED57_2_buffer[clk] != PRED57_2_buffer[!clk]) ||(PRED57_3_buffer[clk] != PRED57_3_buffer[!clk]) ||(PRED57_4_buffer[clk] != PRED57_4_buffer[!clk]) ||(PRED57_5_buffer[clk] != PRED57_5_buffer[!clk]) ||(PRED57_6_buffer[clk] != PRED57_6_buffer[!clk]) ||(PRED57_7_buffer[clk] != PRED57_7_buffer[!clk]) ||(PRED57_8_buffer[clk] != PRED57_8_buffer[!clk]) ||(PRED57_9_buffer[clk] != PRED57_9_buffer[!clk]) ||(PRED57_10_buffer[clk] != PRED57_10_buffer[!clk]) ||(PRED57_11_buffer[clk] != PRED57_11_buffer[!clk]) ||(PRED57_12_buffer[clk] != PRED57_12_buffer[!clk]) ||(PRED57_13_buffer[clk] != PRED57_13_buffer[!clk]) ||(PRED57_14_buffer[clk] != PRED57_14_buffer[!clk]) ||(PRED57_15_buffer[clk] != PRED57_15_buffer[!clk]) ||(PRED57_16_buffer[clk] != PRED57_16_buffer[!clk]) ||(PRED57_17_buffer[clk] != PRED57_17_buffer[!clk]) ||(PRED57_18_buffer[clk] != PRED57_18_buffer[!clk]) ||(PRED57_19_buffer[clk] != PRED57_19_buffer[!clk]) ||(PRED57_20_buffer[clk] != PRED57_20_buffer[!clk]) ||(PRED57_21_buffer[clk] != PRED57_21_buffer[!clk]) ||(PRED57_22_buffer[clk] != PRED57_22_buffer[!clk]) ||(PRED57_23_buffer[clk] != PRED57_23_buffer[!clk]) ||(PRED57_24_buffer[clk] != PRED57_24_buffer[!clk]) ||(PRED57_25_buffer[clk] != PRED57_25_buffer[!clk]) ||(PRED57_26_buffer[clk] != PRED57_26_buffer[!clk]) ||(PRED57_27_buffer[clk] != PRED57_27_buffer[!clk]) ||(PRED57_28_buffer[clk] != PRED57_28_buffer[!clk]) ||(PRED57_29_buffer[clk] != PRED57_29_buffer[!clk]) ||(PRED57_30_buffer[clk] != PRED57_30_buffer[!clk]) ||(PRED57_31_buffer[clk] != PRED57_31_buffer[!clk]) ) begin
      warp1_sig = 1'b1;
    end else begin
      warp1_sig = 1'b0;
    end

    if ((PRED2_0_buffer[clk] != PRED2_0_buffer[!clk]) ||(PRED2_1_buffer[clk] != PRED2_1_buffer[!clk]) ||(PRED2_2_buffer[clk] != PRED2_2_buffer[!clk]) ||(PRED2_3_buffer[clk] != PRED2_3_buffer[!clk]) ||(PRED2_4_buffer[clk] != PRED2_4_buffer[!clk]) ||(PRED2_5_buffer[clk] != PRED2_5_buffer[!clk]) ||(PRED2_6_buffer[clk] != PRED2_6_buffer[!clk]) ||(PRED2_7_buffer[clk] != PRED2_7_buffer[!clk]) ||(PRED2_8_buffer[clk] != PRED2_8_buffer[!clk]) ||(PRED2_9_buffer[clk] != PRED2_9_buffer[!clk]) ||(PRED2_10_buffer[clk] != PRED2_10_buffer[!clk]) ||(PRED2_11_buffer[clk] != PRED2_11_buffer[!clk]) ||(PRED2_12_buffer[clk] != PRED2_12_buffer[!clk]) ||(PRED2_13_buffer[clk] != PRED2_13_buffer[!clk]) ||(PRED2_14_buffer[clk] != PRED2_14_buffer[!clk]) ||(PRED2_15_buffer[clk] != PRED2_15_buffer[!clk]) ||(PRED2_16_buffer[clk] != PRED2_16_buffer[!clk]) ||(PRED2_17_buffer[clk] != PRED2_17_buffer[!clk]) ||(PRED2_18_buffer[clk] != PRED2_18_buffer[!clk]) ||(PRED2_19_buffer[clk] != PRED2_19_buffer[!clk]) ||(PRED2_20_buffer[clk] != PRED2_20_buffer[!clk]) ||(PRED2_21_buffer[clk] != PRED2_21_buffer[!clk]) ||(PRED2_22_buffer[clk] != PRED2_22_buffer[!clk]) ||(PRED2_23_buffer[clk] != PRED2_23_buffer[!clk]) ||(PRED2_24_buffer[clk] != PRED2_24_buffer[!clk]) ||(PRED2_25_buffer[clk] != PRED2_25_buffer[!clk]) ||(PRED2_26_buffer[clk] != PRED2_26_buffer[!clk]) ||(PRED2_27_buffer[clk] != PRED2_27_buffer[!clk]) ||(PRED2_28_buffer[clk] != PRED2_28_buffer[!clk]) ||(PRED2_29_buffer[clk] != PRED2_29_buffer[!clk]) ||(PRED2_30_buffer[clk] != PRED2_30_buffer[!clk]) ||(PRED2_31_buffer[clk] != PRED2_31_buffer[!clk]) ||(PRED10_0_buffer[clk] != PRED10_0_buffer[!clk]) ||(PRED10_1_buffer[clk] != PRED10_1_buffer[!clk]) ||(PRED10_2_buffer[clk] != PRED10_2_buffer[!clk]) ||(PRED10_3_buffer[clk] != PRED10_3_buffer[!clk]) ||(PRED10_4_buffer[clk] != PRED10_4_buffer[!clk]) ||(PRED10_5_buffer[clk] != PRED10_5_buffer[!clk]) ||(PRED10_6_buffer[clk] != PRED10_6_buffer[!clk]) ||(PRED10_7_buffer[clk] != PRED10_7_buffer[!clk]) ||(PRED10_8_buffer[clk] != PRED10_8_buffer[!clk]) ||(PRED10_9_buffer[clk] != PRED10_9_buffer[!clk]) ||(PRED10_10_buffer[clk] != PRED10_10_buffer[!clk]) ||(PRED10_11_buffer[clk] != PRED10_11_buffer[!clk]) ||(PRED10_12_buffer[clk] != PRED10_12_buffer[!clk]) ||(PRED10_13_buffer[clk] != PRED10_13_buffer[!clk]) ||(PRED10_14_buffer[clk] != PRED10_14_buffer[!clk]) ||(PRED10_15_buffer[clk] != PRED10_15_buffer[!clk]) ||(PRED10_16_buffer[clk] != PRED10_16_buffer[!clk]) ||(PRED10_17_buffer[clk] != PRED10_17_buffer[!clk]) ||(PRED10_18_buffer[clk] != PRED10_18_buffer[!clk]) ||(PRED10_19_buffer[clk] != PRED10_19_buffer[!clk]) ||(PRED10_20_buffer[clk] != PRED10_20_buffer[!clk]) ||(PRED10_21_buffer[clk] != PRED10_21_buffer[!clk]) ||(PRED10_22_buffer[clk] != PRED10_22_buffer[!clk]) ||(PRED10_23_buffer[clk] != PRED10_23_buffer[!clk]) ||(PRED10_24_buffer[clk] != PRED10_24_buffer[!clk]) ||(PRED10_25_buffer[clk] != PRED10_25_buffer[!clk]) ||(PRED10_26_buffer[clk] != PRED10_26_buffer[!clk]) ||(PRED10_27_buffer[clk] != PRED10_27_buffer[!clk]) ||(PRED10_28_buffer[clk] != PRED10_28_buffer[!clk]) ||(PRED10_29_buffer[clk] != PRED10_29_buffer[!clk]) ||(PRED10_30_buffer[clk] != PRED10_30_buffer[!clk]) ||(PRED10_31_buffer[clk] != PRED10_31_buffer[!clk]) ||(PRED18_0_buffer[clk] != PRED18_0_buffer[!clk]) ||(PRED18_1_buffer[clk] != PRED18_1_buffer[!clk]) ||(PRED18_2_buffer[clk] != PRED18_2_buffer[!clk]) ||(PRED18_3_buffer[clk] != PRED18_3_buffer[!clk]) ||(PRED18_4_buffer[clk] != PRED18_4_buffer[!clk]) ||(PRED18_5_buffer[clk] != PRED18_5_buffer[!clk]) ||(PRED18_6_buffer[clk] != PRED18_6_buffer[!clk]) ||(PRED18_7_buffer[clk] != PRED18_7_buffer[!clk]) ||(PRED18_8_buffer[clk] != PRED18_8_buffer[!clk]) ||(PRED18_9_buffer[clk] != PRED18_9_buffer[!clk]) ||(PRED18_10_buffer[clk] != PRED18_10_buffer[!clk]) ||(PRED18_11_buffer[clk] != PRED18_11_buffer[!clk]) ||(PRED18_12_buffer[clk] != PRED18_12_buffer[!clk]) ||(PRED18_13_buffer[clk] != PRED18_13_buffer[!clk]) ||(PRED18_14_buffer[clk] != PRED18_14_buffer[!clk]) ||(PRED18_15_buffer[clk] != PRED18_15_buffer[!clk]) ||(PRED18_16_buffer[clk] != PRED18_16_buffer[!clk]) ||(PRED18_17_buffer[clk] != PRED18_17_buffer[!clk]) ||(PRED18_18_buffer[clk] != PRED18_18_buffer[!clk]) ||(PRED18_19_buffer[clk] != PRED18_19_buffer[!clk]) ||(PRED18_20_buffer[clk] != PRED18_20_buffer[!clk]) ||(PRED18_21_buffer[clk] != PRED18_21_buffer[!clk]) ||(PRED18_22_buffer[clk] != PRED18_22_buffer[!clk]) ||(PRED18_23_buffer[clk] != PRED18_23_buffer[!clk]) ||(PRED18_24_buffer[clk] != PRED18_24_buffer[!clk]) ||(PRED18_25_buffer[clk] != PRED18_25_buffer[!clk]) ||(PRED18_26_buffer[clk] != PRED18_26_buffer[!clk]) ||(PRED18_27_buffer[clk] != PRED18_27_buffer[!clk]) ||(PRED18_28_buffer[clk] != PRED18_28_buffer[!clk]) ||(PRED18_29_buffer[clk] != PRED18_29_buffer[!clk]) ||(PRED18_30_buffer[clk] != PRED18_30_buffer[!clk]) ||(PRED18_31_buffer[clk] != PRED18_31_buffer[!clk]) ||(PRED26_0_buffer[clk] != PRED26_0_buffer[!clk]) ||(PRED26_1_buffer[clk] != PRED26_1_buffer[!clk]) ||(PRED26_2_buffer[clk] != PRED26_2_buffer[!clk]) ||(PRED26_3_buffer[clk] != PRED26_3_buffer[!clk]) ||(PRED26_4_buffer[clk] != PRED26_4_buffer[!clk]) ||(PRED26_5_buffer[clk] != PRED26_5_buffer[!clk]) ||(PRED26_6_buffer[clk] != PRED26_6_buffer[!clk]) ||(PRED26_7_buffer[clk] != PRED26_7_buffer[!clk]) ||(PRED26_8_buffer[clk] != PRED26_8_buffer[!clk]) ||(PRED26_9_buffer[clk] != PRED26_9_buffer[!clk]) ||(PRED26_10_buffer[clk] != PRED26_10_buffer[!clk]) ||(PRED26_11_buffer[clk] != PRED26_11_buffer[!clk]) ||(PRED26_12_buffer[clk] != PRED26_12_buffer[!clk]) ||(PRED26_13_buffer[clk] != PRED26_13_buffer[!clk]) ||(PRED26_14_buffer[clk] != PRED26_14_buffer[!clk]) ||(PRED26_15_buffer[clk] != PRED26_15_buffer[!clk]) ||(PRED26_16_buffer[clk] != PRED26_16_buffer[!clk]) ||(PRED26_17_buffer[clk] != PRED26_17_buffer[!clk]) ||(PRED26_18_buffer[clk] != PRED26_18_buffer[!clk]) ||(PRED26_19_buffer[clk] != PRED26_19_buffer[!clk]) ||(PRED26_20_buffer[clk] != PRED26_20_buffer[!clk]) ||(PRED26_21_buffer[clk] != PRED26_21_buffer[!clk]) ||(PRED26_22_buffer[clk] != PRED26_22_buffer[!clk]) ||(PRED26_23_buffer[clk] != PRED26_23_buffer[!clk]) ||(PRED26_24_buffer[clk] != PRED26_24_buffer[!clk]) ||(PRED26_25_buffer[clk] != PRED26_25_buffer[!clk]) ||(PRED26_26_buffer[clk] != PRED26_26_buffer[!clk]) ||(PRED26_27_buffer[clk] != PRED26_27_buffer[!clk]) ||(PRED26_28_buffer[clk] != PRED26_28_buffer[!clk]) ||(PRED26_29_buffer[clk] != PRED26_29_buffer[!clk]) ||(PRED26_30_buffer[clk] != PRED26_30_buffer[!clk]) ||(PRED26_31_buffer[clk] != PRED26_31_buffer[!clk]) ||(PRED34_0_buffer[clk] != PRED34_0_buffer[!clk]) ||(PRED34_1_buffer[clk] != PRED34_1_buffer[!clk]) ||(PRED34_2_buffer[clk] != PRED34_2_buffer[!clk]) ||(PRED34_3_buffer[clk] != PRED34_3_buffer[!clk]) ||(PRED34_4_buffer[clk] != PRED34_4_buffer[!clk]) ||(PRED34_5_buffer[clk] != PRED34_5_buffer[!clk]) ||(PRED34_6_buffer[clk] != PRED34_6_buffer[!clk]) ||(PRED34_7_buffer[clk] != PRED34_7_buffer[!clk]) ||(PRED34_8_buffer[clk] != PRED34_8_buffer[!clk]) ||(PRED34_9_buffer[clk] != PRED34_9_buffer[!clk]) ||(PRED34_10_buffer[clk] != PRED34_10_buffer[!clk]) ||(PRED34_11_buffer[clk] != PRED34_11_buffer[!clk]) ||(PRED34_12_buffer[clk] != PRED34_12_buffer[!clk]) ||(PRED34_13_buffer[clk] != PRED34_13_buffer[!clk]) ||(PRED34_14_buffer[clk] != PRED34_14_buffer[!clk]) ||(PRED34_15_buffer[clk] != PRED34_15_buffer[!clk]) ||(PRED34_16_buffer[clk] != PRED34_16_buffer[!clk]) ||(PRED34_17_buffer[clk] != PRED34_17_buffer[!clk]) ||(PRED34_18_buffer[clk] != PRED34_18_buffer[!clk]) ||(PRED34_19_buffer[clk] != PRED34_19_buffer[!clk]) ||(PRED34_20_buffer[clk] != PRED34_20_buffer[!clk]) ||(PRED34_21_buffer[clk] != PRED34_21_buffer[!clk]) ||(PRED34_22_buffer[clk] != PRED34_22_buffer[!clk]) ||(PRED34_23_buffer[clk] != PRED34_23_buffer[!clk]) ||(PRED34_24_buffer[clk] != PRED34_24_buffer[!clk]) ||(PRED34_25_buffer[clk] != PRED34_25_buffer[!clk]) ||(PRED34_26_buffer[clk] != PRED34_26_buffer[!clk]) ||(PRED34_27_buffer[clk] != PRED34_27_buffer[!clk]) ||(PRED34_28_buffer[clk] != PRED34_28_buffer[!clk]) ||(PRED34_29_buffer[clk] != PRED34_29_buffer[!clk]) ||(PRED34_30_buffer[clk] != PRED34_30_buffer[!clk]) ||(PRED34_31_buffer[clk] != PRED34_31_buffer[!clk]) ||(PRED42_0_buffer[clk] != PRED42_0_buffer[!clk]) ||(PRED42_1_buffer[clk] != PRED42_1_buffer[!clk]) ||(PRED42_2_buffer[clk] != PRED42_2_buffer[!clk]) ||(PRED42_3_buffer[clk] != PRED42_3_buffer[!clk]) ||(PRED42_4_buffer[clk] != PRED42_4_buffer[!clk]) ||(PRED42_5_buffer[clk] != PRED42_5_buffer[!clk]) ||(PRED42_6_buffer[clk] != PRED42_6_buffer[!clk]) ||(PRED42_7_buffer[clk] != PRED42_7_buffer[!clk]) ||(PRED42_8_buffer[clk] != PRED42_8_buffer[!clk]) ||(PRED42_9_buffer[clk] != PRED42_9_buffer[!clk]) ||(PRED42_10_buffer[clk] != PRED42_10_buffer[!clk]) ||(PRED42_11_buffer[clk] != PRED42_11_buffer[!clk]) ||(PRED42_12_buffer[clk] != PRED42_12_buffer[!clk]) ||(PRED42_13_buffer[clk] != PRED42_13_buffer[!clk]) ||(PRED42_14_buffer[clk] != PRED42_14_buffer[!clk]) ||(PRED42_15_buffer[clk] != PRED42_15_buffer[!clk]) ||(PRED42_16_buffer[clk] != PRED42_16_buffer[!clk]) ||(PRED42_17_buffer[clk] != PRED42_17_buffer[!clk]) ||(PRED42_18_buffer[clk] != PRED42_18_buffer[!clk]) ||(PRED42_19_buffer[clk] != PRED42_19_buffer[!clk]) ||(PRED42_20_buffer[clk] != PRED42_20_buffer[!clk]) ||(PRED42_21_buffer[clk] != PRED42_21_buffer[!clk]) ||(PRED42_22_buffer[clk] != PRED42_22_buffer[!clk]) ||(PRED42_23_buffer[clk] != PRED42_23_buffer[!clk]) ||(PRED42_24_buffer[clk] != PRED42_24_buffer[!clk]) ||(PRED42_25_buffer[clk] != PRED42_25_buffer[!clk]) ||(PRED42_26_buffer[clk] != PRED42_26_buffer[!clk]) ||(PRED42_27_buffer[clk] != PRED42_27_buffer[!clk]) ||(PRED42_28_buffer[clk] != PRED42_28_buffer[!clk]) ||(PRED42_29_buffer[clk] != PRED42_29_buffer[!clk]) ||(PRED42_30_buffer[clk] != PRED42_30_buffer[!clk]) ||(PRED42_31_buffer[clk] != PRED42_31_buffer[!clk]) ||(PRED50_0_buffer[clk] != PRED50_0_buffer[!clk]) ||(PRED50_1_buffer[clk] != PRED50_1_buffer[!clk]) ||(PRED50_2_buffer[clk] != PRED50_2_buffer[!clk]) ||(PRED50_3_buffer[clk] != PRED50_3_buffer[!clk]) ||(PRED50_4_buffer[clk] != PRED50_4_buffer[!clk]) ||(PRED50_5_buffer[clk] != PRED50_5_buffer[!clk]) ||(PRED50_6_buffer[clk] != PRED50_6_buffer[!clk]) ||(PRED50_7_buffer[clk] != PRED50_7_buffer[!clk]) ||(PRED50_8_buffer[clk] != PRED50_8_buffer[!clk]) ||(PRED50_9_buffer[clk] != PRED50_9_buffer[!clk]) ||(PRED50_10_buffer[clk] != PRED50_10_buffer[!clk]) ||(PRED50_11_buffer[clk] != PRED50_11_buffer[!clk]) ||(PRED50_12_buffer[clk] != PRED50_12_buffer[!clk]) ||(PRED50_13_buffer[clk] != PRED50_13_buffer[!clk]) ||(PRED50_14_buffer[clk] != PRED50_14_buffer[!clk]) ||(PRED50_15_buffer[clk] != PRED50_15_buffer[!clk]) ||(PRED50_16_buffer[clk] != PRED50_16_buffer[!clk]) ||(PRED50_17_buffer[clk] != PRED50_17_buffer[!clk]) ||(PRED50_18_buffer[clk] != PRED50_18_buffer[!clk]) ||(PRED50_19_buffer[clk] != PRED50_19_buffer[!clk]) ||(PRED50_20_buffer[clk] != PRED50_20_buffer[!clk]) ||(PRED50_21_buffer[clk] != PRED50_21_buffer[!clk]) ||(PRED50_22_buffer[clk] != PRED50_22_buffer[!clk]) ||(PRED50_23_buffer[clk] != PRED50_23_buffer[!clk]) ||(PRED50_24_buffer[clk] != PRED50_24_buffer[!clk]) ||(PRED50_25_buffer[clk] != PRED50_25_buffer[!clk]) ||(PRED50_26_buffer[clk] != PRED50_26_buffer[!clk]) ||(PRED50_27_buffer[clk] != PRED50_27_buffer[!clk]) ||(PRED50_28_buffer[clk] != PRED50_28_buffer[!clk]) ||(PRED50_29_buffer[clk] != PRED50_29_buffer[!clk]) ||(PRED50_30_buffer[clk] != PRED50_30_buffer[!clk]) ||(PRED50_31_buffer[clk] != PRED50_31_buffer[!clk]) ||(PRED58_0_buffer[clk] != PRED58_0_buffer[!clk]) ||(PRED58_1_buffer[clk] != PRED58_1_buffer[!clk]) ||(PRED58_2_buffer[clk] != PRED58_2_buffer[!clk]) ||(PRED58_3_buffer[clk] != PRED58_3_buffer[!clk]) ||(PRED58_4_buffer[clk] != PRED58_4_buffer[!clk]) ||(PRED58_5_buffer[clk] != PRED58_5_buffer[!clk]) ||(PRED58_6_buffer[clk] != PRED58_6_buffer[!clk]) ||(PRED58_7_buffer[clk] != PRED58_7_buffer[!clk]) ||(PRED58_8_buffer[clk] != PRED58_8_buffer[!clk]) ||(PRED58_9_buffer[clk] != PRED58_9_buffer[!clk]) ||(PRED58_10_buffer[clk] != PRED58_10_buffer[!clk]) ||(PRED58_11_buffer[clk] != PRED58_11_buffer[!clk]) ||(PRED58_12_buffer[clk] != PRED58_12_buffer[!clk]) ||(PRED58_13_buffer[clk] != PRED58_13_buffer[!clk]) ||(PRED58_14_buffer[clk] != PRED58_14_buffer[!clk]) ||(PRED58_15_buffer[clk] != PRED58_15_buffer[!clk]) ||(PRED58_16_buffer[clk] != PRED58_16_buffer[!clk]) ||(PRED58_17_buffer[clk] != PRED58_17_buffer[!clk]) ||(PRED58_18_buffer[clk] != PRED58_18_buffer[!clk]) ||(PRED58_19_buffer[clk] != PRED58_19_buffer[!clk]) ||(PRED58_20_buffer[clk] != PRED58_20_buffer[!clk]) ||(PRED58_21_buffer[clk] != PRED58_21_buffer[!clk]) ||(PRED58_22_buffer[clk] != PRED58_22_buffer[!clk]) ||(PRED58_23_buffer[clk] != PRED58_23_buffer[!clk]) ||(PRED58_24_buffer[clk] != PRED58_24_buffer[!clk]) ||(PRED58_25_buffer[clk] != PRED58_25_buffer[!clk]) ||(PRED58_26_buffer[clk] != PRED58_26_buffer[!clk]) ||(PRED58_27_buffer[clk] != PRED58_27_buffer[!clk]) ||(PRED58_28_buffer[clk] != PRED58_28_buffer[!clk]) ||(PRED58_29_buffer[clk] != PRED58_29_buffer[!clk]) ||(PRED58_30_buffer[clk] != PRED58_30_buffer[!clk]) ||(PRED58_31_buffer[clk] != PRED58_31_buffer[!clk]) ) begin
      warp2_sig = 1'b1;
    end else begin
      warp2_sig = 1'b0;
    end

    if ((PRED3_0_buffer[clk] != PRED3_0_buffer[!clk]) ||(PRED3_1_buffer[clk] != PRED3_1_buffer[!clk]) ||(PRED3_2_buffer[clk] != PRED3_2_buffer[!clk]) ||(PRED3_3_buffer[clk] != PRED3_3_buffer[!clk]) ||(PRED3_4_buffer[clk] != PRED3_4_buffer[!clk]) ||(PRED3_5_buffer[clk] != PRED3_5_buffer[!clk]) ||(PRED3_6_buffer[clk] != PRED3_6_buffer[!clk]) ||(PRED3_7_buffer[clk] != PRED3_7_buffer[!clk]) ||(PRED3_8_buffer[clk] != PRED3_8_buffer[!clk]) ||(PRED3_9_buffer[clk] != PRED3_9_buffer[!clk]) ||(PRED3_10_buffer[clk] != PRED3_10_buffer[!clk]) ||(PRED3_11_buffer[clk] != PRED3_11_buffer[!clk]) ||(PRED3_12_buffer[clk] != PRED3_12_buffer[!clk]) ||(PRED3_13_buffer[clk] != PRED3_13_buffer[!clk]) ||(PRED3_14_buffer[clk] != PRED3_14_buffer[!clk]) ||(PRED3_15_buffer[clk] != PRED3_15_buffer[!clk]) ||(PRED3_16_buffer[clk] != PRED3_16_buffer[!clk]) ||(PRED3_17_buffer[clk] != PRED3_17_buffer[!clk]) ||(PRED3_18_buffer[clk] != PRED3_18_buffer[!clk]) ||(PRED3_19_buffer[clk] != PRED3_19_buffer[!clk]) ||(PRED3_20_buffer[clk] != PRED3_20_buffer[!clk]) ||(PRED3_21_buffer[clk] != PRED3_21_buffer[!clk]) ||(PRED3_22_buffer[clk] != PRED3_22_buffer[!clk]) ||(PRED3_23_buffer[clk] != PRED3_23_buffer[!clk]) ||(PRED3_24_buffer[clk] != PRED3_24_buffer[!clk]) ||(PRED3_25_buffer[clk] != PRED3_25_buffer[!clk]) ||(PRED3_26_buffer[clk] != PRED3_26_buffer[!clk]) ||(PRED3_27_buffer[clk] != PRED3_27_buffer[!clk]) ||(PRED3_28_buffer[clk] != PRED3_28_buffer[!clk]) ||(PRED3_29_buffer[clk] != PRED3_29_buffer[!clk]) ||(PRED3_30_buffer[clk] != PRED3_30_buffer[!clk]) ||(PRED3_31_buffer[clk] != PRED3_31_buffer[!clk]) ||(PRED11_0_buffer[clk] != PRED11_0_buffer[!clk]) ||(PRED11_1_buffer[clk] != PRED11_1_buffer[!clk]) ||(PRED11_2_buffer[clk] != PRED11_2_buffer[!clk]) ||(PRED11_3_buffer[clk] != PRED11_3_buffer[!clk]) ||(PRED11_4_buffer[clk] != PRED11_4_buffer[!clk]) ||(PRED11_5_buffer[clk] != PRED11_5_buffer[!clk]) ||(PRED11_6_buffer[clk] != PRED11_6_buffer[!clk]) ||(PRED11_7_buffer[clk] != PRED11_7_buffer[!clk]) ||(PRED11_8_buffer[clk] != PRED11_8_buffer[!clk]) ||(PRED11_9_buffer[clk] != PRED11_9_buffer[!clk]) ||(PRED11_10_buffer[clk] != PRED11_10_buffer[!clk]) ||(PRED11_11_buffer[clk] != PRED11_11_buffer[!clk]) ||(PRED11_12_buffer[clk] != PRED11_12_buffer[!clk]) ||(PRED11_13_buffer[clk] != PRED11_13_buffer[!clk]) ||(PRED11_14_buffer[clk] != PRED11_14_buffer[!clk]) ||(PRED11_15_buffer[clk] != PRED11_15_buffer[!clk]) ||(PRED11_16_buffer[clk] != PRED11_16_buffer[!clk]) ||(PRED11_17_buffer[clk] != PRED11_17_buffer[!clk]) ||(PRED11_18_buffer[clk] != PRED11_18_buffer[!clk]) ||(PRED11_19_buffer[clk] != PRED11_19_buffer[!clk]) ||(PRED11_20_buffer[clk] != PRED11_20_buffer[!clk]) ||(PRED11_21_buffer[clk] != PRED11_21_buffer[!clk]) ||(PRED11_22_buffer[clk] != PRED11_22_buffer[!clk]) ||(PRED11_23_buffer[clk] != PRED11_23_buffer[!clk]) ||(PRED11_24_buffer[clk] != PRED11_24_buffer[!clk]) ||(PRED11_25_buffer[clk] != PRED11_25_buffer[!clk]) ||(PRED11_26_buffer[clk] != PRED11_26_buffer[!clk]) ||(PRED11_27_buffer[clk] != PRED11_27_buffer[!clk]) ||(PRED11_28_buffer[clk] != PRED11_28_buffer[!clk]) ||(PRED11_29_buffer[clk] != PRED11_29_buffer[!clk]) ||(PRED11_30_buffer[clk] != PRED11_30_buffer[!clk]) ||(PRED11_31_buffer[clk] != PRED11_31_buffer[!clk]) ||(PRED19_0_buffer[clk] != PRED19_0_buffer[!clk]) ||(PRED19_1_buffer[clk] != PRED19_1_buffer[!clk]) ||(PRED19_2_buffer[clk] != PRED19_2_buffer[!clk]) ||(PRED19_3_buffer[clk] != PRED19_3_buffer[!clk]) ||(PRED19_4_buffer[clk] != PRED19_4_buffer[!clk]) ||(PRED19_5_buffer[clk] != PRED19_5_buffer[!clk]) ||(PRED19_6_buffer[clk] != PRED19_6_buffer[!clk]) ||(PRED19_7_buffer[clk] != PRED19_7_buffer[!clk]) ||(PRED19_8_buffer[clk] != PRED19_8_buffer[!clk]) ||(PRED19_9_buffer[clk] != PRED19_9_buffer[!clk]) ||(PRED19_10_buffer[clk] != PRED19_10_buffer[!clk]) ||(PRED19_11_buffer[clk] != PRED19_11_buffer[!clk]) ||(PRED19_12_buffer[clk] != PRED19_12_buffer[!clk]) ||(PRED19_13_buffer[clk] != PRED19_13_buffer[!clk]) ||(PRED19_14_buffer[clk] != PRED19_14_buffer[!clk]) ||(PRED19_15_buffer[clk] != PRED19_15_buffer[!clk]) ||(PRED19_16_buffer[clk] != PRED19_16_buffer[!clk]) ||(PRED19_17_buffer[clk] != PRED19_17_buffer[!clk]) ||(PRED19_18_buffer[clk] != PRED19_18_buffer[!clk]) ||(PRED19_19_buffer[clk] != PRED19_19_buffer[!clk]) ||(PRED19_20_buffer[clk] != PRED19_20_buffer[!clk]) ||(PRED19_21_buffer[clk] != PRED19_21_buffer[!clk]) ||(PRED19_22_buffer[clk] != PRED19_22_buffer[!clk]) ||(PRED19_23_buffer[clk] != PRED19_23_buffer[!clk]) ||(PRED19_24_buffer[clk] != PRED19_24_buffer[!clk]) ||(PRED19_25_buffer[clk] != PRED19_25_buffer[!clk]) ||(PRED19_26_buffer[clk] != PRED19_26_buffer[!clk]) ||(PRED19_27_buffer[clk] != PRED19_27_buffer[!clk]) ||(PRED19_28_buffer[clk] != PRED19_28_buffer[!clk]) ||(PRED19_29_buffer[clk] != PRED19_29_buffer[!clk]) ||(PRED19_30_buffer[clk] != PRED19_30_buffer[!clk]) ||(PRED19_31_buffer[clk] != PRED19_31_buffer[!clk]) ||(PRED27_0_buffer[clk] != PRED27_0_buffer[!clk]) ||(PRED27_1_buffer[clk] != PRED27_1_buffer[!clk]) ||(PRED27_2_buffer[clk] != PRED27_2_buffer[!clk]) ||(PRED27_3_buffer[clk] != PRED27_3_buffer[!clk]) ||(PRED27_4_buffer[clk] != PRED27_4_buffer[!clk]) ||(PRED27_5_buffer[clk] != PRED27_5_buffer[!clk]) ||(PRED27_6_buffer[clk] != PRED27_6_buffer[!clk]) ||(PRED27_7_buffer[clk] != PRED27_7_buffer[!clk]) ||(PRED27_8_buffer[clk] != PRED27_8_buffer[!clk]) ||(PRED27_9_buffer[clk] != PRED27_9_buffer[!clk]) ||(PRED27_10_buffer[clk] != PRED27_10_buffer[!clk]) ||(PRED27_11_buffer[clk] != PRED27_11_buffer[!clk]) ||(PRED27_12_buffer[clk] != PRED27_12_buffer[!clk]) ||(PRED27_13_buffer[clk] != PRED27_13_buffer[!clk]) ||(PRED27_14_buffer[clk] != PRED27_14_buffer[!clk]) ||(PRED27_15_buffer[clk] != PRED27_15_buffer[!clk]) ||(PRED27_16_buffer[clk] != PRED27_16_buffer[!clk]) ||(PRED27_17_buffer[clk] != PRED27_17_buffer[!clk]) ||(PRED27_18_buffer[clk] != PRED27_18_buffer[!clk]) ||(PRED27_19_buffer[clk] != PRED27_19_buffer[!clk]) ||(PRED27_20_buffer[clk] != PRED27_20_buffer[!clk]) ||(PRED27_21_buffer[clk] != PRED27_21_buffer[!clk]) ||(PRED27_22_buffer[clk] != PRED27_22_buffer[!clk]) ||(PRED27_23_buffer[clk] != PRED27_23_buffer[!clk]) ||(PRED27_24_buffer[clk] != PRED27_24_buffer[!clk]) ||(PRED27_25_buffer[clk] != PRED27_25_buffer[!clk]) ||(PRED27_26_buffer[clk] != PRED27_26_buffer[!clk]) ||(PRED27_27_buffer[clk] != PRED27_27_buffer[!clk]) ||(PRED27_28_buffer[clk] != PRED27_28_buffer[!clk]) ||(PRED27_29_buffer[clk] != PRED27_29_buffer[!clk]) ||(PRED27_30_buffer[clk] != PRED27_30_buffer[!clk]) ||(PRED27_31_buffer[clk] != PRED27_31_buffer[!clk]) ||(PRED35_0_buffer[clk] != PRED35_0_buffer[!clk]) ||(PRED35_1_buffer[clk] != PRED35_1_buffer[!clk]) ||(PRED35_2_buffer[clk] != PRED35_2_buffer[!clk]) ||(PRED35_3_buffer[clk] != PRED35_3_buffer[!clk]) ||(PRED35_4_buffer[clk] != PRED35_4_buffer[!clk]) ||(PRED35_5_buffer[clk] != PRED35_5_buffer[!clk]) ||(PRED35_6_buffer[clk] != PRED35_6_buffer[!clk]) ||(PRED35_7_buffer[clk] != PRED35_7_buffer[!clk]) ||(PRED35_8_buffer[clk] != PRED35_8_buffer[!clk]) ||(PRED35_9_buffer[clk] != PRED35_9_buffer[!clk]) ||(PRED35_10_buffer[clk] != PRED35_10_buffer[!clk]) ||(PRED35_11_buffer[clk] != PRED35_11_buffer[!clk]) ||(PRED35_12_buffer[clk] != PRED35_12_buffer[!clk]) ||(PRED35_13_buffer[clk] != PRED35_13_buffer[!clk]) ||(PRED35_14_buffer[clk] != PRED35_14_buffer[!clk]) ||(PRED35_15_buffer[clk] != PRED35_15_buffer[!clk]) ||(PRED35_16_buffer[clk] != PRED35_16_buffer[!clk]) ||(PRED35_17_buffer[clk] != PRED35_17_buffer[!clk]) ||(PRED35_18_buffer[clk] != PRED35_18_buffer[!clk]) ||(PRED35_19_buffer[clk] != PRED35_19_buffer[!clk]) ||(PRED35_20_buffer[clk] != PRED35_20_buffer[!clk]) ||(PRED35_21_buffer[clk] != PRED35_21_buffer[!clk]) ||(PRED35_22_buffer[clk] != PRED35_22_buffer[!clk]) ||(PRED35_23_buffer[clk] != PRED35_23_buffer[!clk]) ||(PRED35_24_buffer[clk] != PRED35_24_buffer[!clk]) ||(PRED35_25_buffer[clk] != PRED35_25_buffer[!clk]) ||(PRED35_26_buffer[clk] != PRED35_26_buffer[!clk]) ||(PRED35_27_buffer[clk] != PRED35_27_buffer[!clk]) ||(PRED35_28_buffer[clk] != PRED35_28_buffer[!clk]) ||(PRED35_29_buffer[clk] != PRED35_29_buffer[!clk]) ||(PRED35_30_buffer[clk] != PRED35_30_buffer[!clk]) ||(PRED35_31_buffer[clk] != PRED35_31_buffer[!clk]) ||(PRED43_0_buffer[clk] != PRED43_0_buffer[!clk]) ||(PRED43_1_buffer[clk] != PRED43_1_buffer[!clk]) ||(PRED43_2_buffer[clk] != PRED43_2_buffer[!clk]) ||(PRED43_3_buffer[clk] != PRED43_3_buffer[!clk]) ||(PRED43_4_buffer[clk] != PRED43_4_buffer[!clk]) ||(PRED43_5_buffer[clk] != PRED43_5_buffer[!clk]) ||(PRED43_6_buffer[clk] != PRED43_6_buffer[!clk]) ||(PRED43_7_buffer[clk] != PRED43_7_buffer[!clk]) ||(PRED43_8_buffer[clk] != PRED43_8_buffer[!clk]) ||(PRED43_9_buffer[clk] != PRED43_9_buffer[!clk]) ||(PRED43_10_buffer[clk] != PRED43_10_buffer[!clk]) ||(PRED43_11_buffer[clk] != PRED43_11_buffer[!clk]) ||(PRED43_12_buffer[clk] != PRED43_12_buffer[!clk]) ||(PRED43_13_buffer[clk] != PRED43_13_buffer[!clk]) ||(PRED43_14_buffer[clk] != PRED43_14_buffer[!clk]) ||(PRED43_15_buffer[clk] != PRED43_15_buffer[!clk]) ||(PRED43_16_buffer[clk] != PRED43_16_buffer[!clk]) ||(PRED43_17_buffer[clk] != PRED43_17_buffer[!clk]) ||(PRED43_18_buffer[clk] != PRED43_18_buffer[!clk]) ||(PRED43_19_buffer[clk] != PRED43_19_buffer[!clk]) ||(PRED43_20_buffer[clk] != PRED43_20_buffer[!clk]) ||(PRED43_21_buffer[clk] != PRED43_21_buffer[!clk]) ||(PRED43_22_buffer[clk] != PRED43_22_buffer[!clk]) ||(PRED43_23_buffer[clk] != PRED43_23_buffer[!clk]) ||(PRED43_24_buffer[clk] != PRED43_24_buffer[!clk]) ||(PRED43_25_buffer[clk] != PRED43_25_buffer[!clk]) ||(PRED43_26_buffer[clk] != PRED43_26_buffer[!clk]) ||(PRED43_27_buffer[clk] != PRED43_27_buffer[!clk]) ||(PRED43_28_buffer[clk] != PRED43_28_buffer[!clk]) ||(PRED43_29_buffer[clk] != PRED43_29_buffer[!clk]) ||(PRED43_30_buffer[clk] != PRED43_30_buffer[!clk]) ||(PRED43_31_buffer[clk] != PRED43_31_buffer[!clk]) ||(PRED51_0_buffer[clk] != PRED51_0_buffer[!clk]) ||(PRED51_1_buffer[clk] != PRED51_1_buffer[!clk]) ||(PRED51_2_buffer[clk] != PRED51_2_buffer[!clk]) ||(PRED51_3_buffer[clk] != PRED51_3_buffer[!clk]) ||(PRED51_4_buffer[clk] != PRED51_4_buffer[!clk]) ||(PRED51_5_buffer[clk] != PRED51_5_buffer[!clk]) ||(PRED51_6_buffer[clk] != PRED51_6_buffer[!clk]) ||(PRED51_7_buffer[clk] != PRED51_7_buffer[!clk]) ||(PRED51_8_buffer[clk] != PRED51_8_buffer[!clk]) ||(PRED51_9_buffer[clk] != PRED51_9_buffer[!clk]) ||(PRED51_10_buffer[clk] != PRED51_10_buffer[!clk]) ||(PRED51_11_buffer[clk] != PRED51_11_buffer[!clk]) ||(PRED51_12_buffer[clk] != PRED51_12_buffer[!clk]) ||(PRED51_13_buffer[clk] != PRED51_13_buffer[!clk]) ||(PRED51_14_buffer[clk] != PRED51_14_buffer[!clk]) ||(PRED51_15_buffer[clk] != PRED51_15_buffer[!clk]) ||(PRED51_16_buffer[clk] != PRED51_16_buffer[!clk]) ||(PRED51_17_buffer[clk] != PRED51_17_buffer[!clk]) ||(PRED51_18_buffer[clk] != PRED51_18_buffer[!clk]) ||(PRED51_19_buffer[clk] != PRED51_19_buffer[!clk]) ||(PRED51_20_buffer[clk] != PRED51_20_buffer[!clk]) ||(PRED51_21_buffer[clk] != PRED51_21_buffer[!clk]) ||(PRED51_22_buffer[clk] != PRED51_22_buffer[!clk]) ||(PRED51_23_buffer[clk] != PRED51_23_buffer[!clk]) ||(PRED51_24_buffer[clk] != PRED51_24_buffer[!clk]) ||(PRED51_25_buffer[clk] != PRED51_25_buffer[!clk]) ||(PRED51_26_buffer[clk] != PRED51_26_buffer[!clk]) ||(PRED51_27_buffer[clk] != PRED51_27_buffer[!clk]) ||(PRED51_28_buffer[clk] != PRED51_28_buffer[!clk]) ||(PRED51_29_buffer[clk] != PRED51_29_buffer[!clk]) ||(PRED51_30_buffer[clk] != PRED51_30_buffer[!clk]) ||(PRED51_31_buffer[clk] != PRED51_31_buffer[!clk]) ||(PRED59_0_buffer[clk] != PRED59_0_buffer[!clk]) ||(PRED59_1_buffer[clk] != PRED59_1_buffer[!clk]) ||(PRED59_2_buffer[clk] != PRED59_2_buffer[!clk]) ||(PRED59_3_buffer[clk] != PRED59_3_buffer[!clk]) ||(PRED59_4_buffer[clk] != PRED59_4_buffer[!clk]) ||(PRED59_5_buffer[clk] != PRED59_5_buffer[!clk]) ||(PRED59_6_buffer[clk] != PRED59_6_buffer[!clk]) ||(PRED59_7_buffer[clk] != PRED59_7_buffer[!clk]) ||(PRED59_8_buffer[clk] != PRED59_8_buffer[!clk]) ||(PRED59_9_buffer[clk] != PRED59_9_buffer[!clk]) ||(PRED59_10_buffer[clk] != PRED59_10_buffer[!clk]) ||(PRED59_11_buffer[clk] != PRED59_11_buffer[!clk]) ||(PRED59_12_buffer[clk] != PRED59_12_buffer[!clk]) ||(PRED59_13_buffer[clk] != PRED59_13_buffer[!clk]) ||(PRED59_14_buffer[clk] != PRED59_14_buffer[!clk]) ||(PRED59_15_buffer[clk] != PRED59_15_buffer[!clk]) ||(PRED59_16_buffer[clk] != PRED59_16_buffer[!clk]) ||(PRED59_17_buffer[clk] != PRED59_17_buffer[!clk]) ||(PRED59_18_buffer[clk] != PRED59_18_buffer[!clk]) ||(PRED59_19_buffer[clk] != PRED59_19_buffer[!clk]) ||(PRED59_20_buffer[clk] != PRED59_20_buffer[!clk]) ||(PRED59_21_buffer[clk] != PRED59_21_buffer[!clk]) ||(PRED59_22_buffer[clk] != PRED59_22_buffer[!clk]) ||(PRED59_23_buffer[clk] != PRED59_23_buffer[!clk]) ||(PRED59_24_buffer[clk] != PRED59_24_buffer[!clk]) ||(PRED59_25_buffer[clk] != PRED59_25_buffer[!clk]) ||(PRED59_26_buffer[clk] != PRED59_26_buffer[!clk]) ||(PRED59_27_buffer[clk] != PRED59_27_buffer[!clk]) ||(PRED59_28_buffer[clk] != PRED59_28_buffer[!clk]) ||(PRED59_29_buffer[clk] != PRED59_29_buffer[!clk]) ||(PRED59_30_buffer[clk] != PRED59_30_buffer[!clk]) ||(PRED59_31_buffer[clk] != PRED59_31_buffer[!clk]) ) begin
      warp3_sig = 1'b1;
    end else begin
      warp3_sig = 1'b0;
    end

    if ((PRED4_0_buffer[clk] != PRED4_0_buffer[!clk]) ||(PRED4_1_buffer[clk] != PRED4_1_buffer[!clk]) ||(PRED4_2_buffer[clk] != PRED4_2_buffer[!clk]) ||(PRED4_3_buffer[clk] != PRED4_3_buffer[!clk]) ||(PRED4_4_buffer[clk] != PRED4_4_buffer[!clk]) ||(PRED4_5_buffer[clk] != PRED4_5_buffer[!clk]) ||(PRED4_6_buffer[clk] != PRED4_6_buffer[!clk]) ||(PRED4_7_buffer[clk] != PRED4_7_buffer[!clk]) ||(PRED4_8_buffer[clk] != PRED4_8_buffer[!clk]) ||(PRED4_9_buffer[clk] != PRED4_9_buffer[!clk]) ||(PRED4_10_buffer[clk] != PRED4_10_buffer[!clk]) ||(PRED4_11_buffer[clk] != PRED4_11_buffer[!clk]) ||(PRED4_12_buffer[clk] != PRED4_12_buffer[!clk]) ||(PRED4_13_buffer[clk] != PRED4_13_buffer[!clk]) ||(PRED4_14_buffer[clk] != PRED4_14_buffer[!clk]) ||(PRED4_15_buffer[clk] != PRED4_15_buffer[!clk]) ||(PRED4_16_buffer[clk] != PRED4_16_buffer[!clk]) ||(PRED4_17_buffer[clk] != PRED4_17_buffer[!clk]) ||(PRED4_18_buffer[clk] != PRED4_18_buffer[!clk]) ||(PRED4_19_buffer[clk] != PRED4_19_buffer[!clk]) ||(PRED4_20_buffer[clk] != PRED4_20_buffer[!clk]) ||(PRED4_21_buffer[clk] != PRED4_21_buffer[!clk]) ||(PRED4_22_buffer[clk] != PRED4_22_buffer[!clk]) ||(PRED4_23_buffer[clk] != PRED4_23_buffer[!clk]) ||(PRED4_24_buffer[clk] != PRED4_24_buffer[!clk]) ||(PRED4_25_buffer[clk] != PRED4_25_buffer[!clk]) ||(PRED4_26_buffer[clk] != PRED4_26_buffer[!clk]) ||(PRED4_27_buffer[clk] != PRED4_27_buffer[!clk]) ||(PRED4_28_buffer[clk] != PRED4_28_buffer[!clk]) ||(PRED4_29_buffer[clk] != PRED4_29_buffer[!clk]) ||(PRED4_30_buffer[clk] != PRED4_30_buffer[!clk]) ||(PRED4_31_buffer[clk] != PRED4_31_buffer[!clk]) ||(PRED12_0_buffer[clk] != PRED12_0_buffer[!clk]) ||(PRED12_1_buffer[clk] != PRED12_1_buffer[!clk]) ||(PRED12_2_buffer[clk] != PRED12_2_buffer[!clk]) ||(PRED12_3_buffer[clk] != PRED12_3_buffer[!clk]) ||(PRED12_4_buffer[clk] != PRED12_4_buffer[!clk]) ||(PRED12_5_buffer[clk] != PRED12_5_buffer[!clk]) ||(PRED12_6_buffer[clk] != PRED12_6_buffer[!clk]) ||(PRED12_7_buffer[clk] != PRED12_7_buffer[!clk]) ||(PRED12_8_buffer[clk] != PRED12_8_buffer[!clk]) ||(PRED12_9_buffer[clk] != PRED12_9_buffer[!clk]) ||(PRED12_10_buffer[clk] != PRED12_10_buffer[!clk]) ||(PRED12_11_buffer[clk] != PRED12_11_buffer[!clk]) ||(PRED12_12_buffer[clk] != PRED12_12_buffer[!clk]) ||(PRED12_13_buffer[clk] != PRED12_13_buffer[!clk]) ||(PRED12_14_buffer[clk] != PRED12_14_buffer[!clk]) ||(PRED12_15_buffer[clk] != PRED12_15_buffer[!clk]) ||(PRED12_16_buffer[clk] != PRED12_16_buffer[!clk]) ||(PRED12_17_buffer[clk] != PRED12_17_buffer[!clk]) ||(PRED12_18_buffer[clk] != PRED12_18_buffer[!clk]) ||(PRED12_19_buffer[clk] != PRED12_19_buffer[!clk]) ||(PRED12_20_buffer[clk] != PRED12_20_buffer[!clk]) ||(PRED12_21_buffer[clk] != PRED12_21_buffer[!clk]) ||(PRED12_22_buffer[clk] != PRED12_22_buffer[!clk]) ||(PRED12_23_buffer[clk] != PRED12_23_buffer[!clk]) ||(PRED12_24_buffer[clk] != PRED12_24_buffer[!clk]) ||(PRED12_25_buffer[clk] != PRED12_25_buffer[!clk]) ||(PRED12_26_buffer[clk] != PRED12_26_buffer[!clk]) ||(PRED12_27_buffer[clk] != PRED12_27_buffer[!clk]) ||(PRED12_28_buffer[clk] != PRED12_28_buffer[!clk]) ||(PRED12_29_buffer[clk] != PRED12_29_buffer[!clk]) ||(PRED12_30_buffer[clk] != PRED12_30_buffer[!clk]) ||(PRED12_31_buffer[clk] != PRED12_31_buffer[!clk]) ||(PRED20_0_buffer[clk] != PRED20_0_buffer[!clk]) ||(PRED20_1_buffer[clk] != PRED20_1_buffer[!clk]) ||(PRED20_2_buffer[clk] != PRED20_2_buffer[!clk]) ||(PRED20_3_buffer[clk] != PRED20_3_buffer[!clk]) ||(PRED20_4_buffer[clk] != PRED20_4_buffer[!clk]) ||(PRED20_5_buffer[clk] != PRED20_5_buffer[!clk]) ||(PRED20_6_buffer[clk] != PRED20_6_buffer[!clk]) ||(PRED20_7_buffer[clk] != PRED20_7_buffer[!clk]) ||(PRED20_8_buffer[clk] != PRED20_8_buffer[!clk]) ||(PRED20_9_buffer[clk] != PRED20_9_buffer[!clk]) ||(PRED20_10_buffer[clk] != PRED20_10_buffer[!clk]) ||(PRED20_11_buffer[clk] != PRED20_11_buffer[!clk]) ||(PRED20_12_buffer[clk] != PRED20_12_buffer[!clk]) ||(PRED20_13_buffer[clk] != PRED20_13_buffer[!clk]) ||(PRED20_14_buffer[clk] != PRED20_14_buffer[!clk]) ||(PRED20_15_buffer[clk] != PRED20_15_buffer[!clk]) ||(PRED20_16_buffer[clk] != PRED20_16_buffer[!clk]) ||(PRED20_17_buffer[clk] != PRED20_17_buffer[!clk]) ||(PRED20_18_buffer[clk] != PRED20_18_buffer[!clk]) ||(PRED20_19_buffer[clk] != PRED20_19_buffer[!clk]) ||(PRED20_20_buffer[clk] != PRED20_20_buffer[!clk]) ||(PRED20_21_buffer[clk] != PRED20_21_buffer[!clk]) ||(PRED20_22_buffer[clk] != PRED20_22_buffer[!clk]) ||(PRED20_23_buffer[clk] != PRED20_23_buffer[!clk]) ||(PRED20_24_buffer[clk] != PRED20_24_buffer[!clk]) ||(PRED20_25_buffer[clk] != PRED20_25_buffer[!clk]) ||(PRED20_26_buffer[clk] != PRED20_26_buffer[!clk]) ||(PRED20_27_buffer[clk] != PRED20_27_buffer[!clk]) ||(PRED20_28_buffer[clk] != PRED20_28_buffer[!clk]) ||(PRED20_29_buffer[clk] != PRED20_29_buffer[!clk]) ||(PRED20_30_buffer[clk] != PRED20_30_buffer[!clk]) ||(PRED20_31_buffer[clk] != PRED20_31_buffer[!clk]) ||(PRED28_0_buffer[clk] != PRED28_0_buffer[!clk]) ||(PRED28_1_buffer[clk] != PRED28_1_buffer[!clk]) ||(PRED28_2_buffer[clk] != PRED28_2_buffer[!clk]) ||(PRED28_3_buffer[clk] != PRED28_3_buffer[!clk]) ||(PRED28_4_buffer[clk] != PRED28_4_buffer[!clk]) ||(PRED28_5_buffer[clk] != PRED28_5_buffer[!clk]) ||(PRED28_6_buffer[clk] != PRED28_6_buffer[!clk]) ||(PRED28_7_buffer[clk] != PRED28_7_buffer[!clk]) ||(PRED28_8_buffer[clk] != PRED28_8_buffer[!clk]) ||(PRED28_9_buffer[clk] != PRED28_9_buffer[!clk]) ||(PRED28_10_buffer[clk] != PRED28_10_buffer[!clk]) ||(PRED28_11_buffer[clk] != PRED28_11_buffer[!clk]) ||(PRED28_12_buffer[clk] != PRED28_12_buffer[!clk]) ||(PRED28_13_buffer[clk] != PRED28_13_buffer[!clk]) ||(PRED28_14_buffer[clk] != PRED28_14_buffer[!clk]) ||(PRED28_15_buffer[clk] != PRED28_15_buffer[!clk]) ||(PRED28_16_buffer[clk] != PRED28_16_buffer[!clk]) ||(PRED28_17_buffer[clk] != PRED28_17_buffer[!clk]) ||(PRED28_18_buffer[clk] != PRED28_18_buffer[!clk]) ||(PRED28_19_buffer[clk] != PRED28_19_buffer[!clk]) ||(PRED28_20_buffer[clk] != PRED28_20_buffer[!clk]) ||(PRED28_21_buffer[clk] != PRED28_21_buffer[!clk]) ||(PRED28_22_buffer[clk] != PRED28_22_buffer[!clk]) ||(PRED28_23_buffer[clk] != PRED28_23_buffer[!clk]) ||(PRED28_24_buffer[clk] != PRED28_24_buffer[!clk]) ||(PRED28_25_buffer[clk] != PRED28_25_buffer[!clk]) ||(PRED28_26_buffer[clk] != PRED28_26_buffer[!clk]) ||(PRED28_27_buffer[clk] != PRED28_27_buffer[!clk]) ||(PRED28_28_buffer[clk] != PRED28_28_buffer[!clk]) ||(PRED28_29_buffer[clk] != PRED28_29_buffer[!clk]) ||(PRED28_30_buffer[clk] != PRED28_30_buffer[!clk]) ||(PRED28_31_buffer[clk] != PRED28_31_buffer[!clk]) ||(PRED36_0_buffer[clk] != PRED36_0_buffer[!clk]) ||(PRED36_1_buffer[clk] != PRED36_1_buffer[!clk]) ||(PRED36_2_buffer[clk] != PRED36_2_buffer[!clk]) ||(PRED36_3_buffer[clk] != PRED36_3_buffer[!clk]) ||(PRED36_4_buffer[clk] != PRED36_4_buffer[!clk]) ||(PRED36_5_buffer[clk] != PRED36_5_buffer[!clk]) ||(PRED36_6_buffer[clk] != PRED36_6_buffer[!clk]) ||(PRED36_7_buffer[clk] != PRED36_7_buffer[!clk]) ||(PRED36_8_buffer[clk] != PRED36_8_buffer[!clk]) ||(PRED36_9_buffer[clk] != PRED36_9_buffer[!clk]) ||(PRED36_10_buffer[clk] != PRED36_10_buffer[!clk]) ||(PRED36_11_buffer[clk] != PRED36_11_buffer[!clk]) ||(PRED36_12_buffer[clk] != PRED36_12_buffer[!clk]) ||(PRED36_13_buffer[clk] != PRED36_13_buffer[!clk]) ||(PRED36_14_buffer[clk] != PRED36_14_buffer[!clk]) ||(PRED36_15_buffer[clk] != PRED36_15_buffer[!clk]) ||(PRED36_16_buffer[clk] != PRED36_16_buffer[!clk]) ||(PRED36_17_buffer[clk] != PRED36_17_buffer[!clk]) ||(PRED36_18_buffer[clk] != PRED36_18_buffer[!clk]) ||(PRED36_19_buffer[clk] != PRED36_19_buffer[!clk]) ||(PRED36_20_buffer[clk] != PRED36_20_buffer[!clk]) ||(PRED36_21_buffer[clk] != PRED36_21_buffer[!clk]) ||(PRED36_22_buffer[clk] != PRED36_22_buffer[!clk]) ||(PRED36_23_buffer[clk] != PRED36_23_buffer[!clk]) ||(PRED36_24_buffer[clk] != PRED36_24_buffer[!clk]) ||(PRED36_25_buffer[clk] != PRED36_25_buffer[!clk]) ||(PRED36_26_buffer[clk] != PRED36_26_buffer[!clk]) ||(PRED36_27_buffer[clk] != PRED36_27_buffer[!clk]) ||(PRED36_28_buffer[clk] != PRED36_28_buffer[!clk]) ||(PRED36_29_buffer[clk] != PRED36_29_buffer[!clk]) ||(PRED36_30_buffer[clk] != PRED36_30_buffer[!clk]) ||(PRED36_31_buffer[clk] != PRED36_31_buffer[!clk]) ||(PRED44_0_buffer[clk] != PRED44_0_buffer[!clk]) ||(PRED44_1_buffer[clk] != PRED44_1_buffer[!clk]) ||(PRED44_2_buffer[clk] != PRED44_2_buffer[!clk]) ||(PRED44_3_buffer[clk] != PRED44_3_buffer[!clk]) ||(PRED44_4_buffer[clk] != PRED44_4_buffer[!clk]) ||(PRED44_5_buffer[clk] != PRED44_5_buffer[!clk]) ||(PRED44_6_buffer[clk] != PRED44_6_buffer[!clk]) ||(PRED44_7_buffer[clk] != PRED44_7_buffer[!clk]) ||(PRED44_8_buffer[clk] != PRED44_8_buffer[!clk]) ||(PRED44_9_buffer[clk] != PRED44_9_buffer[!clk]) ||(PRED44_10_buffer[clk] != PRED44_10_buffer[!clk]) ||(PRED44_11_buffer[clk] != PRED44_11_buffer[!clk]) ||(PRED44_12_buffer[clk] != PRED44_12_buffer[!clk]) ||(PRED44_13_buffer[clk] != PRED44_13_buffer[!clk]) ||(PRED44_14_buffer[clk] != PRED44_14_buffer[!clk]) ||(PRED44_15_buffer[clk] != PRED44_15_buffer[!clk]) ||(PRED44_16_buffer[clk] != PRED44_16_buffer[!clk]) ||(PRED44_17_buffer[clk] != PRED44_17_buffer[!clk]) ||(PRED44_18_buffer[clk] != PRED44_18_buffer[!clk]) ||(PRED44_19_buffer[clk] != PRED44_19_buffer[!clk]) ||(PRED44_20_buffer[clk] != PRED44_20_buffer[!clk]) ||(PRED44_21_buffer[clk] != PRED44_21_buffer[!clk]) ||(PRED44_22_buffer[clk] != PRED44_22_buffer[!clk]) ||(PRED44_23_buffer[clk] != PRED44_23_buffer[!clk]) ||(PRED44_24_buffer[clk] != PRED44_24_buffer[!clk]) ||(PRED44_25_buffer[clk] != PRED44_25_buffer[!clk]) ||(PRED44_26_buffer[clk] != PRED44_26_buffer[!clk]) ||(PRED44_27_buffer[clk] != PRED44_27_buffer[!clk]) ||(PRED44_28_buffer[clk] != PRED44_28_buffer[!clk]) ||(PRED44_29_buffer[clk] != PRED44_29_buffer[!clk]) ||(PRED44_30_buffer[clk] != PRED44_30_buffer[!clk]) ||(PRED44_31_buffer[clk] != PRED44_31_buffer[!clk]) ||(PRED52_0_buffer[clk] != PRED52_0_buffer[!clk]) ||(PRED52_1_buffer[clk] != PRED52_1_buffer[!clk]) ||(PRED52_2_buffer[clk] != PRED52_2_buffer[!clk]) ||(PRED52_3_buffer[clk] != PRED52_3_buffer[!clk]) ||(PRED52_4_buffer[clk] != PRED52_4_buffer[!clk]) ||(PRED52_5_buffer[clk] != PRED52_5_buffer[!clk]) ||(PRED52_6_buffer[clk] != PRED52_6_buffer[!clk]) ||(PRED52_7_buffer[clk] != PRED52_7_buffer[!clk]) ||(PRED52_8_buffer[clk] != PRED52_8_buffer[!clk]) ||(PRED52_9_buffer[clk] != PRED52_9_buffer[!clk]) ||(PRED52_10_buffer[clk] != PRED52_10_buffer[!clk]) ||(PRED52_11_buffer[clk] != PRED52_11_buffer[!clk]) ||(PRED52_12_buffer[clk] != PRED52_12_buffer[!clk]) ||(PRED52_13_buffer[clk] != PRED52_13_buffer[!clk]) ||(PRED52_14_buffer[clk] != PRED52_14_buffer[!clk]) ||(PRED52_15_buffer[clk] != PRED52_15_buffer[!clk]) ||(PRED52_16_buffer[clk] != PRED52_16_buffer[!clk]) ||(PRED52_17_buffer[clk] != PRED52_17_buffer[!clk]) ||(PRED52_18_buffer[clk] != PRED52_18_buffer[!clk]) ||(PRED52_19_buffer[clk] != PRED52_19_buffer[!clk]) ||(PRED52_20_buffer[clk] != PRED52_20_buffer[!clk]) ||(PRED52_21_buffer[clk] != PRED52_21_buffer[!clk]) ||(PRED52_22_buffer[clk] != PRED52_22_buffer[!clk]) ||(PRED52_23_buffer[clk] != PRED52_23_buffer[!clk]) ||(PRED52_24_buffer[clk] != PRED52_24_buffer[!clk]) ||(PRED52_25_buffer[clk] != PRED52_25_buffer[!clk]) ||(PRED52_26_buffer[clk] != PRED52_26_buffer[!clk]) ||(PRED52_27_buffer[clk] != PRED52_27_buffer[!clk]) ||(PRED52_28_buffer[clk] != PRED52_28_buffer[!clk]) ||(PRED52_29_buffer[clk] != PRED52_29_buffer[!clk]) ||(PRED52_30_buffer[clk] != PRED52_30_buffer[!clk]) ||(PRED52_31_buffer[clk] != PRED52_31_buffer[!clk]) ||(PRED60_0_buffer[clk] != PRED60_0_buffer[!clk]) ||(PRED60_1_buffer[clk] != PRED60_1_buffer[!clk]) ||(PRED60_2_buffer[clk] != PRED60_2_buffer[!clk]) ||(PRED60_3_buffer[clk] != PRED60_3_buffer[!clk]) ||(PRED60_4_buffer[clk] != PRED60_4_buffer[!clk]) ||(PRED60_5_buffer[clk] != PRED60_5_buffer[!clk]) ||(PRED60_6_buffer[clk] != PRED60_6_buffer[!clk]) ||(PRED60_7_buffer[clk] != PRED60_7_buffer[!clk]) ||(PRED60_8_buffer[clk] != PRED60_8_buffer[!clk]) ||(PRED60_9_buffer[clk] != PRED60_9_buffer[!clk]) ||(PRED60_10_buffer[clk] != PRED60_10_buffer[!clk]) ||(PRED60_11_buffer[clk] != PRED60_11_buffer[!clk]) ||(PRED60_12_buffer[clk] != PRED60_12_buffer[!clk]) ||(PRED60_13_buffer[clk] != PRED60_13_buffer[!clk]) ||(PRED60_14_buffer[clk] != PRED60_14_buffer[!clk]) ||(PRED60_15_buffer[clk] != PRED60_15_buffer[!clk]) ||(PRED60_16_buffer[clk] != PRED60_16_buffer[!clk]) ||(PRED60_17_buffer[clk] != PRED60_17_buffer[!clk]) ||(PRED60_18_buffer[clk] != PRED60_18_buffer[!clk]) ||(PRED60_19_buffer[clk] != PRED60_19_buffer[!clk]) ||(PRED60_20_buffer[clk] != PRED60_20_buffer[!clk]) ||(PRED60_21_buffer[clk] != PRED60_21_buffer[!clk]) ||(PRED60_22_buffer[clk] != PRED60_22_buffer[!clk]) ||(PRED60_23_buffer[clk] != PRED60_23_buffer[!clk]) ||(PRED60_24_buffer[clk] != PRED60_24_buffer[!clk]) ||(PRED60_25_buffer[clk] != PRED60_25_buffer[!clk]) ||(PRED60_26_buffer[clk] != PRED60_26_buffer[!clk]) ||(PRED60_27_buffer[clk] != PRED60_27_buffer[!clk]) ||(PRED60_28_buffer[clk] != PRED60_28_buffer[!clk]) ||(PRED60_29_buffer[clk] != PRED60_29_buffer[!clk]) ||(PRED60_30_buffer[clk] != PRED60_30_buffer[!clk]) ||(PRED60_31_buffer[clk] != PRED60_31_buffer[!clk]) ) begin
      warp4_sig = 1'b1;
    end else begin
      warp4_sig = 1'b0;
    end

    if ((PRED5_0_buffer[clk] != PRED5_0_buffer[!clk]) ||(PRED5_1_buffer[clk] != PRED5_1_buffer[!clk]) ||(PRED5_2_buffer[clk] != PRED5_2_buffer[!clk]) ||(PRED5_3_buffer[clk] != PRED5_3_buffer[!clk]) ||(PRED5_4_buffer[clk] != PRED5_4_buffer[!clk]) ||(PRED5_5_buffer[clk] != PRED5_5_buffer[!clk]) ||(PRED5_6_buffer[clk] != PRED5_6_buffer[!clk]) ||(PRED5_7_buffer[clk] != PRED5_7_buffer[!clk]) ||(PRED5_8_buffer[clk] != PRED5_8_buffer[!clk]) ||(PRED5_9_buffer[clk] != PRED5_9_buffer[!clk]) ||(PRED5_10_buffer[clk] != PRED5_10_buffer[!clk]) ||(PRED5_11_buffer[clk] != PRED5_11_buffer[!clk]) ||(PRED5_12_buffer[clk] != PRED5_12_buffer[!clk]) ||(PRED5_13_buffer[clk] != PRED5_13_buffer[!clk]) ||(PRED5_14_buffer[clk] != PRED5_14_buffer[!clk]) ||(PRED5_15_buffer[clk] != PRED5_15_buffer[!clk]) ||(PRED5_16_buffer[clk] != PRED5_16_buffer[!clk]) ||(PRED5_17_buffer[clk] != PRED5_17_buffer[!clk]) ||(PRED5_18_buffer[clk] != PRED5_18_buffer[!clk]) ||(PRED5_19_buffer[clk] != PRED5_19_buffer[!clk]) ||(PRED5_20_buffer[clk] != PRED5_20_buffer[!clk]) ||(PRED5_21_buffer[clk] != PRED5_21_buffer[!clk]) ||(PRED5_22_buffer[clk] != PRED5_22_buffer[!clk]) ||(PRED5_23_buffer[clk] != PRED5_23_buffer[!clk]) ||(PRED5_24_buffer[clk] != PRED5_24_buffer[!clk]) ||(PRED5_25_buffer[clk] != PRED5_25_buffer[!clk]) ||(PRED5_26_buffer[clk] != PRED5_26_buffer[!clk]) ||(PRED5_27_buffer[clk] != PRED5_27_buffer[!clk]) ||(PRED5_28_buffer[clk] != PRED5_28_buffer[!clk]) ||(PRED5_29_buffer[clk] != PRED5_29_buffer[!clk]) ||(PRED5_30_buffer[clk] != PRED5_30_buffer[!clk]) ||(PRED5_31_buffer[clk] != PRED5_31_buffer[!clk]) ||(PRED13_0_buffer[clk] != PRED13_0_buffer[!clk]) ||(PRED13_1_buffer[clk] != PRED13_1_buffer[!clk]) ||(PRED13_2_buffer[clk] != PRED13_2_buffer[!clk]) ||(PRED13_3_buffer[clk] != PRED13_3_buffer[!clk]) ||(PRED13_4_buffer[clk] != PRED13_4_buffer[!clk]) ||(PRED13_5_buffer[clk] != PRED13_5_buffer[!clk]) ||(PRED13_6_buffer[clk] != PRED13_6_buffer[!clk]) ||(PRED13_7_buffer[clk] != PRED13_7_buffer[!clk]) ||(PRED13_8_buffer[clk] != PRED13_8_buffer[!clk]) ||(PRED13_9_buffer[clk] != PRED13_9_buffer[!clk]) ||(PRED13_10_buffer[clk] != PRED13_10_buffer[!clk]) ||(PRED13_11_buffer[clk] != PRED13_11_buffer[!clk]) ||(PRED13_12_buffer[clk] != PRED13_12_buffer[!clk]) ||(PRED13_13_buffer[clk] != PRED13_13_buffer[!clk]) ||(PRED13_14_buffer[clk] != PRED13_14_buffer[!clk]) ||(PRED13_15_buffer[clk] != PRED13_15_buffer[!clk]) ||(PRED13_16_buffer[clk] != PRED13_16_buffer[!clk]) ||(PRED13_17_buffer[clk] != PRED13_17_buffer[!clk]) ||(PRED13_18_buffer[clk] != PRED13_18_buffer[!clk]) ||(PRED13_19_buffer[clk] != PRED13_19_buffer[!clk]) ||(PRED13_20_buffer[clk] != PRED13_20_buffer[!clk]) ||(PRED13_21_buffer[clk] != PRED13_21_buffer[!clk]) ||(PRED13_22_buffer[clk] != PRED13_22_buffer[!clk]) ||(PRED13_23_buffer[clk] != PRED13_23_buffer[!clk]) ||(PRED13_24_buffer[clk] != PRED13_24_buffer[!clk]) ||(PRED13_25_buffer[clk] != PRED13_25_buffer[!clk]) ||(PRED13_26_buffer[clk] != PRED13_26_buffer[!clk]) ||(PRED13_27_buffer[clk] != PRED13_27_buffer[!clk]) ||(PRED13_28_buffer[clk] != PRED13_28_buffer[!clk]) ||(PRED13_29_buffer[clk] != PRED13_29_buffer[!clk]) ||(PRED13_30_buffer[clk] != PRED13_30_buffer[!clk]) ||(PRED13_31_buffer[clk] != PRED13_31_buffer[!clk]) ||(PRED21_0_buffer[clk] != PRED21_0_buffer[!clk]) ||(PRED21_1_buffer[clk] != PRED21_1_buffer[!clk]) ||(PRED21_2_buffer[clk] != PRED21_2_buffer[!clk]) ||(PRED21_3_buffer[clk] != PRED21_3_buffer[!clk]) ||(PRED21_4_buffer[clk] != PRED21_4_buffer[!clk]) ||(PRED21_5_buffer[clk] != PRED21_5_buffer[!clk]) ||(PRED21_6_buffer[clk] != PRED21_6_buffer[!clk]) ||(PRED21_7_buffer[clk] != PRED21_7_buffer[!clk]) ||(PRED21_8_buffer[clk] != PRED21_8_buffer[!clk]) ||(PRED21_9_buffer[clk] != PRED21_9_buffer[!clk]) ||(PRED21_10_buffer[clk] != PRED21_10_buffer[!clk]) ||(PRED21_11_buffer[clk] != PRED21_11_buffer[!clk]) ||(PRED21_12_buffer[clk] != PRED21_12_buffer[!clk]) ||(PRED21_13_buffer[clk] != PRED21_13_buffer[!clk]) ||(PRED21_14_buffer[clk] != PRED21_14_buffer[!clk]) ||(PRED21_15_buffer[clk] != PRED21_15_buffer[!clk]) ||(PRED21_16_buffer[clk] != PRED21_16_buffer[!clk]) ||(PRED21_17_buffer[clk] != PRED21_17_buffer[!clk]) ||(PRED21_18_buffer[clk] != PRED21_18_buffer[!clk]) ||(PRED21_19_buffer[clk] != PRED21_19_buffer[!clk]) ||(PRED21_20_buffer[clk] != PRED21_20_buffer[!clk]) ||(PRED21_21_buffer[clk] != PRED21_21_buffer[!clk]) ||(PRED21_22_buffer[clk] != PRED21_22_buffer[!clk]) ||(PRED21_23_buffer[clk] != PRED21_23_buffer[!clk]) ||(PRED21_24_buffer[clk] != PRED21_24_buffer[!clk]) ||(PRED21_25_buffer[clk] != PRED21_25_buffer[!clk]) ||(PRED21_26_buffer[clk] != PRED21_26_buffer[!clk]) ||(PRED21_27_buffer[clk] != PRED21_27_buffer[!clk]) ||(PRED21_28_buffer[clk] != PRED21_28_buffer[!clk]) ||(PRED21_29_buffer[clk] != PRED21_29_buffer[!clk]) ||(PRED21_30_buffer[clk] != PRED21_30_buffer[!clk]) ||(PRED21_31_buffer[clk] != PRED21_31_buffer[!clk]) ||(PRED29_0_buffer[clk] != PRED29_0_buffer[!clk]) ||(PRED29_1_buffer[clk] != PRED29_1_buffer[!clk]) ||(PRED29_2_buffer[clk] != PRED29_2_buffer[!clk]) ||(PRED29_3_buffer[clk] != PRED29_3_buffer[!clk]) ||(PRED29_4_buffer[clk] != PRED29_4_buffer[!clk]) ||(PRED29_5_buffer[clk] != PRED29_5_buffer[!clk]) ||(PRED29_6_buffer[clk] != PRED29_6_buffer[!clk]) ||(PRED29_7_buffer[clk] != PRED29_7_buffer[!clk]) ||(PRED29_8_buffer[clk] != PRED29_8_buffer[!clk]) ||(PRED29_9_buffer[clk] != PRED29_9_buffer[!clk]) ||(PRED29_10_buffer[clk] != PRED29_10_buffer[!clk]) ||(PRED29_11_buffer[clk] != PRED29_11_buffer[!clk]) ||(PRED29_12_buffer[clk] != PRED29_12_buffer[!clk]) ||(PRED29_13_buffer[clk] != PRED29_13_buffer[!clk]) ||(PRED29_14_buffer[clk] != PRED29_14_buffer[!clk]) ||(PRED29_15_buffer[clk] != PRED29_15_buffer[!clk]) ||(PRED29_16_buffer[clk] != PRED29_16_buffer[!clk]) ||(PRED29_17_buffer[clk] != PRED29_17_buffer[!clk]) ||(PRED29_18_buffer[clk] != PRED29_18_buffer[!clk]) ||(PRED29_19_buffer[clk] != PRED29_19_buffer[!clk]) ||(PRED29_20_buffer[clk] != PRED29_20_buffer[!clk]) ||(PRED29_21_buffer[clk] != PRED29_21_buffer[!clk]) ||(PRED29_22_buffer[clk] != PRED29_22_buffer[!clk]) ||(PRED29_23_buffer[clk] != PRED29_23_buffer[!clk]) ||(PRED29_24_buffer[clk] != PRED29_24_buffer[!clk]) ||(PRED29_25_buffer[clk] != PRED29_25_buffer[!clk]) ||(PRED29_26_buffer[clk] != PRED29_26_buffer[!clk]) ||(PRED29_27_buffer[clk] != PRED29_27_buffer[!clk]) ||(PRED29_28_buffer[clk] != PRED29_28_buffer[!clk]) ||(PRED29_29_buffer[clk] != PRED29_29_buffer[!clk]) ||(PRED29_30_buffer[clk] != PRED29_30_buffer[!clk]) ||(PRED29_31_buffer[clk] != PRED29_31_buffer[!clk]) ||(PRED37_0_buffer[clk] != PRED37_0_buffer[!clk]) ||(PRED37_1_buffer[clk] != PRED37_1_buffer[!clk]) ||(PRED37_2_buffer[clk] != PRED37_2_buffer[!clk]) ||(PRED37_3_buffer[clk] != PRED37_3_buffer[!clk]) ||(PRED37_4_buffer[clk] != PRED37_4_buffer[!clk]) ||(PRED37_5_buffer[clk] != PRED37_5_buffer[!clk]) ||(PRED37_6_buffer[clk] != PRED37_6_buffer[!clk]) ||(PRED37_7_buffer[clk] != PRED37_7_buffer[!clk]) ||(PRED37_8_buffer[clk] != PRED37_8_buffer[!clk]) ||(PRED37_9_buffer[clk] != PRED37_9_buffer[!clk]) ||(PRED37_10_buffer[clk] != PRED37_10_buffer[!clk]) ||(PRED37_11_buffer[clk] != PRED37_11_buffer[!clk]) ||(PRED37_12_buffer[clk] != PRED37_12_buffer[!clk]) ||(PRED37_13_buffer[clk] != PRED37_13_buffer[!clk]) ||(PRED37_14_buffer[clk] != PRED37_14_buffer[!clk]) ||(PRED37_15_buffer[clk] != PRED37_15_buffer[!clk]) ||(PRED37_16_buffer[clk] != PRED37_16_buffer[!clk]) ||(PRED37_17_buffer[clk] != PRED37_17_buffer[!clk]) ||(PRED37_18_buffer[clk] != PRED37_18_buffer[!clk]) ||(PRED37_19_buffer[clk] != PRED37_19_buffer[!clk]) ||(PRED37_20_buffer[clk] != PRED37_20_buffer[!clk]) ||(PRED37_21_buffer[clk] != PRED37_21_buffer[!clk]) ||(PRED37_22_buffer[clk] != PRED37_22_buffer[!clk]) ||(PRED37_23_buffer[clk] != PRED37_23_buffer[!clk]) ||(PRED37_24_buffer[clk] != PRED37_24_buffer[!clk]) ||(PRED37_25_buffer[clk] != PRED37_25_buffer[!clk]) ||(PRED37_26_buffer[clk] != PRED37_26_buffer[!clk]) ||(PRED37_27_buffer[clk] != PRED37_27_buffer[!clk]) ||(PRED37_28_buffer[clk] != PRED37_28_buffer[!clk]) ||(PRED37_29_buffer[clk] != PRED37_29_buffer[!clk]) ||(PRED37_30_buffer[clk] != PRED37_30_buffer[!clk]) ||(PRED37_31_buffer[clk] != PRED37_31_buffer[!clk]) ||(PRED45_0_buffer[clk] != PRED45_0_buffer[!clk]) ||(PRED45_1_buffer[clk] != PRED45_1_buffer[!clk]) ||(PRED45_2_buffer[clk] != PRED45_2_buffer[!clk]) ||(PRED45_3_buffer[clk] != PRED45_3_buffer[!clk]) ||(PRED45_4_buffer[clk] != PRED45_4_buffer[!clk]) ||(PRED45_5_buffer[clk] != PRED45_5_buffer[!clk]) ||(PRED45_6_buffer[clk] != PRED45_6_buffer[!clk]) ||(PRED45_7_buffer[clk] != PRED45_7_buffer[!clk]) ||(PRED45_8_buffer[clk] != PRED45_8_buffer[!clk]) ||(PRED45_9_buffer[clk] != PRED45_9_buffer[!clk]) ||(PRED45_10_buffer[clk] != PRED45_10_buffer[!clk]) ||(PRED45_11_buffer[clk] != PRED45_11_buffer[!clk]) ||(PRED45_12_buffer[clk] != PRED45_12_buffer[!clk]) ||(PRED45_13_buffer[clk] != PRED45_13_buffer[!clk]) ||(PRED45_14_buffer[clk] != PRED45_14_buffer[!clk]) ||(PRED45_15_buffer[clk] != PRED45_15_buffer[!clk]) ||(PRED45_16_buffer[clk] != PRED45_16_buffer[!clk]) ||(PRED45_17_buffer[clk] != PRED45_17_buffer[!clk]) ||(PRED45_18_buffer[clk] != PRED45_18_buffer[!clk]) ||(PRED45_19_buffer[clk] != PRED45_19_buffer[!clk]) ||(PRED45_20_buffer[clk] != PRED45_20_buffer[!clk]) ||(PRED45_21_buffer[clk] != PRED45_21_buffer[!clk]) ||(PRED45_22_buffer[clk] != PRED45_22_buffer[!clk]) ||(PRED45_23_buffer[clk] != PRED45_23_buffer[!clk]) ||(PRED45_24_buffer[clk] != PRED45_24_buffer[!clk]) ||(PRED45_25_buffer[clk] != PRED45_25_buffer[!clk]) ||(PRED45_26_buffer[clk] != PRED45_26_buffer[!clk]) ||(PRED45_27_buffer[clk] != PRED45_27_buffer[!clk]) ||(PRED45_28_buffer[clk] != PRED45_28_buffer[!clk]) ||(PRED45_29_buffer[clk] != PRED45_29_buffer[!clk]) ||(PRED45_30_buffer[clk] != PRED45_30_buffer[!clk]) ||(PRED45_31_buffer[clk] != PRED45_31_buffer[!clk]) ||(PRED53_0_buffer[clk] != PRED53_0_buffer[!clk]) ||(PRED53_1_buffer[clk] != PRED53_1_buffer[!clk]) ||(PRED53_2_buffer[clk] != PRED53_2_buffer[!clk]) ||(PRED53_3_buffer[clk] != PRED53_3_buffer[!clk]) ||(PRED53_4_buffer[clk] != PRED53_4_buffer[!clk]) ||(PRED53_5_buffer[clk] != PRED53_5_buffer[!clk]) ||(PRED53_6_buffer[clk] != PRED53_6_buffer[!clk]) ||(PRED53_7_buffer[clk] != PRED53_7_buffer[!clk]) ||(PRED53_8_buffer[clk] != PRED53_8_buffer[!clk]) ||(PRED53_9_buffer[clk] != PRED53_9_buffer[!clk]) ||(PRED53_10_buffer[clk] != PRED53_10_buffer[!clk]) ||(PRED53_11_buffer[clk] != PRED53_11_buffer[!clk]) ||(PRED53_12_buffer[clk] != PRED53_12_buffer[!clk]) ||(PRED53_13_buffer[clk] != PRED53_13_buffer[!clk]) ||(PRED53_14_buffer[clk] != PRED53_14_buffer[!clk]) ||(PRED53_15_buffer[clk] != PRED53_15_buffer[!clk]) ||(PRED53_16_buffer[clk] != PRED53_16_buffer[!clk]) ||(PRED53_17_buffer[clk] != PRED53_17_buffer[!clk]) ||(PRED53_18_buffer[clk] != PRED53_18_buffer[!clk]) ||(PRED53_19_buffer[clk] != PRED53_19_buffer[!clk]) ||(PRED53_20_buffer[clk] != PRED53_20_buffer[!clk]) ||(PRED53_21_buffer[clk] != PRED53_21_buffer[!clk]) ||(PRED53_22_buffer[clk] != PRED53_22_buffer[!clk]) ||(PRED53_23_buffer[clk] != PRED53_23_buffer[!clk]) ||(PRED53_24_buffer[clk] != PRED53_24_buffer[!clk]) ||(PRED53_25_buffer[clk] != PRED53_25_buffer[!clk]) ||(PRED53_26_buffer[clk] != PRED53_26_buffer[!clk]) ||(PRED53_27_buffer[clk] != PRED53_27_buffer[!clk]) ||(PRED53_28_buffer[clk] != PRED53_28_buffer[!clk]) ||(PRED53_29_buffer[clk] != PRED53_29_buffer[!clk]) ||(PRED53_30_buffer[clk] != PRED53_30_buffer[!clk]) ||(PRED53_31_buffer[clk] != PRED53_31_buffer[!clk]) ||(PRED61_0_buffer[clk] != PRED61_0_buffer[!clk]) ||(PRED61_1_buffer[clk] != PRED61_1_buffer[!clk]) ||(PRED61_2_buffer[clk] != PRED61_2_buffer[!clk]) ||(PRED61_3_buffer[clk] != PRED61_3_buffer[!clk]) ||(PRED61_4_buffer[clk] != PRED61_4_buffer[!clk]) ||(PRED61_5_buffer[clk] != PRED61_5_buffer[!clk]) ||(PRED61_6_buffer[clk] != PRED61_6_buffer[!clk]) ||(PRED61_7_buffer[clk] != PRED61_7_buffer[!clk]) ||(PRED61_8_buffer[clk] != PRED61_8_buffer[!clk]) ||(PRED61_9_buffer[clk] != PRED61_9_buffer[!clk]) ||(PRED61_10_buffer[clk] != PRED61_10_buffer[!clk]) ||(PRED61_11_buffer[clk] != PRED61_11_buffer[!clk]) ||(PRED61_12_buffer[clk] != PRED61_12_buffer[!clk]) ||(PRED61_13_buffer[clk] != PRED61_13_buffer[!clk]) ||(PRED61_14_buffer[clk] != PRED61_14_buffer[!clk]) ||(PRED61_15_buffer[clk] != PRED61_15_buffer[!clk]) ||(PRED61_16_buffer[clk] != PRED61_16_buffer[!clk]) ||(PRED61_17_buffer[clk] != PRED61_17_buffer[!clk]) ||(PRED61_18_buffer[clk] != PRED61_18_buffer[!clk]) ||(PRED61_19_buffer[clk] != PRED61_19_buffer[!clk]) ||(PRED61_20_buffer[clk] != PRED61_20_buffer[!clk]) ||(PRED61_21_buffer[clk] != PRED61_21_buffer[!clk]) ||(PRED61_22_buffer[clk] != PRED61_22_buffer[!clk]) ||(PRED61_23_buffer[clk] != PRED61_23_buffer[!clk]) ||(PRED61_24_buffer[clk] != PRED61_24_buffer[!clk]) ||(PRED61_25_buffer[clk] != PRED61_25_buffer[!clk]) ||(PRED61_26_buffer[clk] != PRED61_26_buffer[!clk]) ||(PRED61_27_buffer[clk] != PRED61_27_buffer[!clk]) ||(PRED61_28_buffer[clk] != PRED61_28_buffer[!clk]) ||(PRED61_29_buffer[clk] != PRED61_29_buffer[!clk]) ||(PRED61_30_buffer[clk] != PRED61_30_buffer[!clk]) ||(PRED61_31_buffer[clk] != PRED61_31_buffer[!clk]) ) begin
      warp5_sig = 1'b1;
    end else begin
      warp5_sig = 1'b0;
    end

    if ((PRED6_0_buffer[clk] != PRED6_0_buffer[!clk]) ||(PRED6_1_buffer[clk] != PRED6_1_buffer[!clk]) ||(PRED6_2_buffer[clk] != PRED6_2_buffer[!clk]) ||(PRED6_3_buffer[clk] != PRED6_3_buffer[!clk]) ||(PRED6_4_buffer[clk] != PRED6_4_buffer[!clk]) ||(PRED6_5_buffer[clk] != PRED6_5_buffer[!clk]) ||(PRED6_6_buffer[clk] != PRED6_6_buffer[!clk]) ||(PRED6_7_buffer[clk] != PRED6_7_buffer[!clk]) ||(PRED6_8_buffer[clk] != PRED6_8_buffer[!clk]) ||(PRED6_9_buffer[clk] != PRED6_9_buffer[!clk]) ||(PRED6_10_buffer[clk] != PRED6_10_buffer[!clk]) ||(PRED6_11_buffer[clk] != PRED6_11_buffer[!clk]) ||(PRED6_12_buffer[clk] != PRED6_12_buffer[!clk]) ||(PRED6_13_buffer[clk] != PRED6_13_buffer[!clk]) ||(PRED6_14_buffer[clk] != PRED6_14_buffer[!clk]) ||(PRED6_15_buffer[clk] != PRED6_15_buffer[!clk]) ||(PRED6_16_buffer[clk] != PRED6_16_buffer[!clk]) ||(PRED6_17_buffer[clk] != PRED6_17_buffer[!clk]) ||(PRED6_18_buffer[clk] != PRED6_18_buffer[!clk]) ||(PRED6_19_buffer[clk] != PRED6_19_buffer[!clk]) ||(PRED6_20_buffer[clk] != PRED6_20_buffer[!clk]) ||(PRED6_21_buffer[clk] != PRED6_21_buffer[!clk]) ||(PRED6_22_buffer[clk] != PRED6_22_buffer[!clk]) ||(PRED6_23_buffer[clk] != PRED6_23_buffer[!clk]) ||(PRED6_24_buffer[clk] != PRED6_24_buffer[!clk]) ||(PRED6_25_buffer[clk] != PRED6_25_buffer[!clk]) ||(PRED6_26_buffer[clk] != PRED6_26_buffer[!clk]) ||(PRED6_27_buffer[clk] != PRED6_27_buffer[!clk]) ||(PRED6_28_buffer[clk] != PRED6_28_buffer[!clk]) ||(PRED6_29_buffer[clk] != PRED6_29_buffer[!clk]) ||(PRED6_30_buffer[clk] != PRED6_30_buffer[!clk]) ||(PRED6_31_buffer[clk] != PRED6_31_buffer[!clk]) ||(PRED14_0_buffer[clk] != PRED14_0_buffer[!clk]) ||(PRED14_1_buffer[clk] != PRED14_1_buffer[!clk]) ||(PRED14_2_buffer[clk] != PRED14_2_buffer[!clk]) ||(PRED14_3_buffer[clk] != PRED14_3_buffer[!clk]) ||(PRED14_4_buffer[clk] != PRED14_4_buffer[!clk]) ||(PRED14_5_buffer[clk] != PRED14_5_buffer[!clk]) ||(PRED14_6_buffer[clk] != PRED14_6_buffer[!clk]) ||(PRED14_7_buffer[clk] != PRED14_7_buffer[!clk]) ||(PRED14_8_buffer[clk] != PRED14_8_buffer[!clk]) ||(PRED14_9_buffer[clk] != PRED14_9_buffer[!clk]) ||(PRED14_10_buffer[clk] != PRED14_10_buffer[!clk]) ||(PRED14_11_buffer[clk] != PRED14_11_buffer[!clk]) ||(PRED14_12_buffer[clk] != PRED14_12_buffer[!clk]) ||(PRED14_13_buffer[clk] != PRED14_13_buffer[!clk]) ||(PRED14_14_buffer[clk] != PRED14_14_buffer[!clk]) ||(PRED14_15_buffer[clk] != PRED14_15_buffer[!clk]) ||(PRED14_16_buffer[clk] != PRED14_16_buffer[!clk]) ||(PRED14_17_buffer[clk] != PRED14_17_buffer[!clk]) ||(PRED14_18_buffer[clk] != PRED14_18_buffer[!clk]) ||(PRED14_19_buffer[clk] != PRED14_19_buffer[!clk]) ||(PRED14_20_buffer[clk] != PRED14_20_buffer[!clk]) ||(PRED14_21_buffer[clk] != PRED14_21_buffer[!clk]) ||(PRED14_22_buffer[clk] != PRED14_22_buffer[!clk]) ||(PRED14_23_buffer[clk] != PRED14_23_buffer[!clk]) ||(PRED14_24_buffer[clk] != PRED14_24_buffer[!clk]) ||(PRED14_25_buffer[clk] != PRED14_25_buffer[!clk]) ||(PRED14_26_buffer[clk] != PRED14_26_buffer[!clk]) ||(PRED14_27_buffer[clk] != PRED14_27_buffer[!clk]) ||(PRED14_28_buffer[clk] != PRED14_28_buffer[!clk]) ||(PRED14_29_buffer[clk] != PRED14_29_buffer[!clk]) ||(PRED14_30_buffer[clk] != PRED14_30_buffer[!clk]) ||(PRED14_31_buffer[clk] != PRED14_31_buffer[!clk]) ||(PRED22_0_buffer[clk] != PRED22_0_buffer[!clk]) ||(PRED22_1_buffer[clk] != PRED22_1_buffer[!clk]) ||(PRED22_2_buffer[clk] != PRED22_2_buffer[!clk]) ||(PRED22_3_buffer[clk] != PRED22_3_buffer[!clk]) ||(PRED22_4_buffer[clk] != PRED22_4_buffer[!clk]) ||(PRED22_5_buffer[clk] != PRED22_5_buffer[!clk]) ||(PRED22_6_buffer[clk] != PRED22_6_buffer[!clk]) ||(PRED22_7_buffer[clk] != PRED22_7_buffer[!clk]) ||(PRED22_8_buffer[clk] != PRED22_8_buffer[!clk]) ||(PRED22_9_buffer[clk] != PRED22_9_buffer[!clk]) ||(PRED22_10_buffer[clk] != PRED22_10_buffer[!clk]) ||(PRED22_11_buffer[clk] != PRED22_11_buffer[!clk]) ||(PRED22_12_buffer[clk] != PRED22_12_buffer[!clk]) ||(PRED22_13_buffer[clk] != PRED22_13_buffer[!clk]) ||(PRED22_14_buffer[clk] != PRED22_14_buffer[!clk]) ||(PRED22_15_buffer[clk] != PRED22_15_buffer[!clk]) ||(PRED22_16_buffer[clk] != PRED22_16_buffer[!clk]) ||(PRED22_17_buffer[clk] != PRED22_17_buffer[!clk]) ||(PRED22_18_buffer[clk] != PRED22_18_buffer[!clk]) ||(PRED22_19_buffer[clk] != PRED22_19_buffer[!clk]) ||(PRED22_20_buffer[clk] != PRED22_20_buffer[!clk]) ||(PRED22_21_buffer[clk] != PRED22_21_buffer[!clk]) ||(PRED22_22_buffer[clk] != PRED22_22_buffer[!clk]) ||(PRED22_23_buffer[clk] != PRED22_23_buffer[!clk]) ||(PRED22_24_buffer[clk] != PRED22_24_buffer[!clk]) ||(PRED22_25_buffer[clk] != PRED22_25_buffer[!clk]) ||(PRED22_26_buffer[clk] != PRED22_26_buffer[!clk]) ||(PRED22_27_buffer[clk] != PRED22_27_buffer[!clk]) ||(PRED22_28_buffer[clk] != PRED22_28_buffer[!clk]) ||(PRED22_29_buffer[clk] != PRED22_29_buffer[!clk]) ||(PRED22_30_buffer[clk] != PRED22_30_buffer[!clk]) ||(PRED22_31_buffer[clk] != PRED22_31_buffer[!clk]) ||(PRED30_0_buffer[clk] != PRED30_0_buffer[!clk]) ||(PRED30_1_buffer[clk] != PRED30_1_buffer[!clk]) ||(PRED30_2_buffer[clk] != PRED30_2_buffer[!clk]) ||(PRED30_3_buffer[clk] != PRED30_3_buffer[!clk]) ||(PRED30_4_buffer[clk] != PRED30_4_buffer[!clk]) ||(PRED30_5_buffer[clk] != PRED30_5_buffer[!clk]) ||(PRED30_6_buffer[clk] != PRED30_6_buffer[!clk]) ||(PRED30_7_buffer[clk] != PRED30_7_buffer[!clk]) ||(PRED30_8_buffer[clk] != PRED30_8_buffer[!clk]) ||(PRED30_9_buffer[clk] != PRED30_9_buffer[!clk]) ||(PRED30_10_buffer[clk] != PRED30_10_buffer[!clk]) ||(PRED30_11_buffer[clk] != PRED30_11_buffer[!clk]) ||(PRED30_12_buffer[clk] != PRED30_12_buffer[!clk]) ||(PRED30_13_buffer[clk] != PRED30_13_buffer[!clk]) ||(PRED30_14_buffer[clk] != PRED30_14_buffer[!clk]) ||(PRED30_15_buffer[clk] != PRED30_15_buffer[!clk]) ||(PRED30_16_buffer[clk] != PRED30_16_buffer[!clk]) ||(PRED30_17_buffer[clk] != PRED30_17_buffer[!clk]) ||(PRED30_18_buffer[clk] != PRED30_18_buffer[!clk]) ||(PRED30_19_buffer[clk] != PRED30_19_buffer[!clk]) ||(PRED30_20_buffer[clk] != PRED30_20_buffer[!clk]) ||(PRED30_21_buffer[clk] != PRED30_21_buffer[!clk]) ||(PRED30_22_buffer[clk] != PRED30_22_buffer[!clk]) ||(PRED30_23_buffer[clk] != PRED30_23_buffer[!clk]) ||(PRED30_24_buffer[clk] != PRED30_24_buffer[!clk]) ||(PRED30_25_buffer[clk] != PRED30_25_buffer[!clk]) ||(PRED30_26_buffer[clk] != PRED30_26_buffer[!clk]) ||(PRED30_27_buffer[clk] != PRED30_27_buffer[!clk]) ||(PRED30_28_buffer[clk] != PRED30_28_buffer[!clk]) ||(PRED30_29_buffer[clk] != PRED30_29_buffer[!clk]) ||(PRED30_30_buffer[clk] != PRED30_30_buffer[!clk]) ||(PRED30_31_buffer[clk] != PRED30_31_buffer[!clk]) ||(PRED38_0_buffer[clk] != PRED38_0_buffer[!clk]) ||(PRED38_1_buffer[clk] != PRED38_1_buffer[!clk]) ||(PRED38_2_buffer[clk] != PRED38_2_buffer[!clk]) ||(PRED38_3_buffer[clk] != PRED38_3_buffer[!clk]) ||(PRED38_4_buffer[clk] != PRED38_4_buffer[!clk]) ||(PRED38_5_buffer[clk] != PRED38_5_buffer[!clk]) ||(PRED38_6_buffer[clk] != PRED38_6_buffer[!clk]) ||(PRED38_7_buffer[clk] != PRED38_7_buffer[!clk]) ||(PRED38_8_buffer[clk] != PRED38_8_buffer[!clk]) ||(PRED38_9_buffer[clk] != PRED38_9_buffer[!clk]) ||(PRED38_10_buffer[clk] != PRED38_10_buffer[!clk]) ||(PRED38_11_buffer[clk] != PRED38_11_buffer[!clk]) ||(PRED38_12_buffer[clk] != PRED38_12_buffer[!clk]) ||(PRED38_13_buffer[clk] != PRED38_13_buffer[!clk]) ||(PRED38_14_buffer[clk] != PRED38_14_buffer[!clk]) ||(PRED38_15_buffer[clk] != PRED38_15_buffer[!clk]) ||(PRED38_16_buffer[clk] != PRED38_16_buffer[!clk]) ||(PRED38_17_buffer[clk] != PRED38_17_buffer[!clk]) ||(PRED38_18_buffer[clk] != PRED38_18_buffer[!clk]) ||(PRED38_19_buffer[clk] != PRED38_19_buffer[!clk]) ||(PRED38_20_buffer[clk] != PRED38_20_buffer[!clk]) ||(PRED38_21_buffer[clk] != PRED38_21_buffer[!clk]) ||(PRED38_22_buffer[clk] != PRED38_22_buffer[!clk]) ||(PRED38_23_buffer[clk] != PRED38_23_buffer[!clk]) ||(PRED38_24_buffer[clk] != PRED38_24_buffer[!clk]) ||(PRED38_25_buffer[clk] != PRED38_25_buffer[!clk]) ||(PRED38_26_buffer[clk] != PRED38_26_buffer[!clk]) ||(PRED38_27_buffer[clk] != PRED38_27_buffer[!clk]) ||(PRED38_28_buffer[clk] != PRED38_28_buffer[!clk]) ||(PRED38_29_buffer[clk] != PRED38_29_buffer[!clk]) ||(PRED38_30_buffer[clk] != PRED38_30_buffer[!clk]) ||(PRED38_31_buffer[clk] != PRED38_31_buffer[!clk]) ||(PRED46_0_buffer[clk] != PRED46_0_buffer[!clk]) ||(PRED46_1_buffer[clk] != PRED46_1_buffer[!clk]) ||(PRED46_2_buffer[clk] != PRED46_2_buffer[!clk]) ||(PRED46_3_buffer[clk] != PRED46_3_buffer[!clk]) ||(PRED46_4_buffer[clk] != PRED46_4_buffer[!clk]) ||(PRED46_5_buffer[clk] != PRED46_5_buffer[!clk]) ||(PRED46_6_buffer[clk] != PRED46_6_buffer[!clk]) ||(PRED46_7_buffer[clk] != PRED46_7_buffer[!clk]) ||(PRED46_8_buffer[clk] != PRED46_8_buffer[!clk]) ||(PRED46_9_buffer[clk] != PRED46_9_buffer[!clk]) ||(PRED46_10_buffer[clk] != PRED46_10_buffer[!clk]) ||(PRED46_11_buffer[clk] != PRED46_11_buffer[!clk]) ||(PRED46_12_buffer[clk] != PRED46_12_buffer[!clk]) ||(PRED46_13_buffer[clk] != PRED46_13_buffer[!clk]) ||(PRED46_14_buffer[clk] != PRED46_14_buffer[!clk]) ||(PRED46_15_buffer[clk] != PRED46_15_buffer[!clk]) ||(PRED46_16_buffer[clk] != PRED46_16_buffer[!clk]) ||(PRED46_17_buffer[clk] != PRED46_17_buffer[!clk]) ||(PRED46_18_buffer[clk] != PRED46_18_buffer[!clk]) ||(PRED46_19_buffer[clk] != PRED46_19_buffer[!clk]) ||(PRED46_20_buffer[clk] != PRED46_20_buffer[!clk]) ||(PRED46_21_buffer[clk] != PRED46_21_buffer[!clk]) ||(PRED46_22_buffer[clk] != PRED46_22_buffer[!clk]) ||(PRED46_23_buffer[clk] != PRED46_23_buffer[!clk]) ||(PRED46_24_buffer[clk] != PRED46_24_buffer[!clk]) ||(PRED46_25_buffer[clk] != PRED46_25_buffer[!clk]) ||(PRED46_26_buffer[clk] != PRED46_26_buffer[!clk]) ||(PRED46_27_buffer[clk] != PRED46_27_buffer[!clk]) ||(PRED46_28_buffer[clk] != PRED46_28_buffer[!clk]) ||(PRED46_29_buffer[clk] != PRED46_29_buffer[!clk]) ||(PRED46_30_buffer[clk] != PRED46_30_buffer[!clk]) ||(PRED46_31_buffer[clk] != PRED46_31_buffer[!clk]) ||(PRED54_0_buffer[clk] != PRED54_0_buffer[!clk]) ||(PRED54_1_buffer[clk] != PRED54_1_buffer[!clk]) ||(PRED54_2_buffer[clk] != PRED54_2_buffer[!clk]) ||(PRED54_3_buffer[clk] != PRED54_3_buffer[!clk]) ||(PRED54_4_buffer[clk] != PRED54_4_buffer[!clk]) ||(PRED54_5_buffer[clk] != PRED54_5_buffer[!clk]) ||(PRED54_6_buffer[clk] != PRED54_6_buffer[!clk]) ||(PRED54_7_buffer[clk] != PRED54_7_buffer[!clk]) ||(PRED54_8_buffer[clk] != PRED54_8_buffer[!clk]) ||(PRED54_9_buffer[clk] != PRED54_9_buffer[!clk]) ||(PRED54_10_buffer[clk] != PRED54_10_buffer[!clk]) ||(PRED54_11_buffer[clk] != PRED54_11_buffer[!clk]) ||(PRED54_12_buffer[clk] != PRED54_12_buffer[!clk]) ||(PRED54_13_buffer[clk] != PRED54_13_buffer[!clk]) ||(PRED54_14_buffer[clk] != PRED54_14_buffer[!clk]) ||(PRED54_15_buffer[clk] != PRED54_15_buffer[!clk]) ||(PRED54_16_buffer[clk] != PRED54_16_buffer[!clk]) ||(PRED54_17_buffer[clk] != PRED54_17_buffer[!clk]) ||(PRED54_18_buffer[clk] != PRED54_18_buffer[!clk]) ||(PRED54_19_buffer[clk] != PRED54_19_buffer[!clk]) ||(PRED54_20_buffer[clk] != PRED54_20_buffer[!clk]) ||(PRED54_21_buffer[clk] != PRED54_21_buffer[!clk]) ||(PRED54_22_buffer[clk] != PRED54_22_buffer[!clk]) ||(PRED54_23_buffer[clk] != PRED54_23_buffer[!clk]) ||(PRED54_24_buffer[clk] != PRED54_24_buffer[!clk]) ||(PRED54_25_buffer[clk] != PRED54_25_buffer[!clk]) ||(PRED54_26_buffer[clk] != PRED54_26_buffer[!clk]) ||(PRED54_27_buffer[clk] != PRED54_27_buffer[!clk]) ||(PRED54_28_buffer[clk] != PRED54_28_buffer[!clk]) ||(PRED54_29_buffer[clk] != PRED54_29_buffer[!clk]) ||(PRED54_30_buffer[clk] != PRED54_30_buffer[!clk]) ||(PRED54_31_buffer[clk] != PRED54_31_buffer[!clk]) ||(PRED62_0_buffer[clk] != PRED62_0_buffer[!clk]) ||(PRED62_1_buffer[clk] != PRED62_1_buffer[!clk]) ||(PRED62_2_buffer[clk] != PRED62_2_buffer[!clk]) ||(PRED62_3_buffer[clk] != PRED62_3_buffer[!clk]) ||(PRED62_4_buffer[clk] != PRED62_4_buffer[!clk]) ||(PRED62_5_buffer[clk] != PRED62_5_buffer[!clk]) ||(PRED62_6_buffer[clk] != PRED62_6_buffer[!clk]) ||(PRED62_7_buffer[clk] != PRED62_7_buffer[!clk]) ||(PRED62_8_buffer[clk] != PRED62_8_buffer[!clk]) ||(PRED62_9_buffer[clk] != PRED62_9_buffer[!clk]) ||(PRED62_10_buffer[clk] != PRED62_10_buffer[!clk]) ||(PRED62_11_buffer[clk] != PRED62_11_buffer[!clk]) ||(PRED62_12_buffer[clk] != PRED62_12_buffer[!clk]) ||(PRED62_13_buffer[clk] != PRED62_13_buffer[!clk]) ||(PRED62_14_buffer[clk] != PRED62_14_buffer[!clk]) ||(PRED62_15_buffer[clk] != PRED62_15_buffer[!clk]) ||(PRED62_16_buffer[clk] != PRED62_16_buffer[!clk]) ||(PRED62_17_buffer[clk] != PRED62_17_buffer[!clk]) ||(PRED62_18_buffer[clk] != PRED62_18_buffer[!clk]) ||(PRED62_19_buffer[clk] != PRED62_19_buffer[!clk]) ||(PRED62_20_buffer[clk] != PRED62_20_buffer[!clk]) ||(PRED62_21_buffer[clk] != PRED62_21_buffer[!clk]) ||(PRED62_22_buffer[clk] != PRED62_22_buffer[!clk]) ||(PRED62_23_buffer[clk] != PRED62_23_buffer[!clk]) ||(PRED62_24_buffer[clk] != PRED62_24_buffer[!clk]) ||(PRED62_25_buffer[clk] != PRED62_25_buffer[!clk]) ||(PRED62_26_buffer[clk] != PRED62_26_buffer[!clk]) ||(PRED62_27_buffer[clk] != PRED62_27_buffer[!clk]) ||(PRED62_28_buffer[clk] != PRED62_28_buffer[!clk]) ||(PRED62_29_buffer[clk] != PRED62_29_buffer[!clk]) ||(PRED62_30_buffer[clk] != PRED62_30_buffer[!clk]) ||(PRED62_31_buffer[clk] != PRED62_31_buffer[!clk]) ) begin
      warp6_sig = 1'b1;
    end else begin
      warp6_sig = 1'b0;
    end

    if ((PRED7_0_buffer[clk] != PRED7_0_buffer[!clk]) ||(PRED7_1_buffer[clk] != PRED7_1_buffer[!clk]) ||(PRED7_2_buffer[clk] != PRED7_2_buffer[!clk]) ||(PRED7_3_buffer[clk] != PRED7_3_buffer[!clk]) ||(PRED7_4_buffer[clk] != PRED7_4_buffer[!clk]) ||(PRED7_5_buffer[clk] != PRED7_5_buffer[!clk]) ||(PRED7_6_buffer[clk] != PRED7_6_buffer[!clk]) ||(PRED7_7_buffer[clk] != PRED7_7_buffer[!clk]) ||(PRED7_8_buffer[clk] != PRED7_8_buffer[!clk]) ||(PRED7_9_buffer[clk] != PRED7_9_buffer[!clk]) ||(PRED7_10_buffer[clk] != PRED7_10_buffer[!clk]) ||(PRED7_11_buffer[clk] != PRED7_11_buffer[!clk]) ||(PRED7_12_buffer[clk] != PRED7_12_buffer[!clk]) ||(PRED7_13_buffer[clk] != PRED7_13_buffer[!clk]) ||(PRED7_14_buffer[clk] != PRED7_14_buffer[!clk]) ||(PRED7_15_buffer[clk] != PRED7_15_buffer[!clk]) ||(PRED7_16_buffer[clk] != PRED7_16_buffer[!clk]) ||(PRED7_17_buffer[clk] != PRED7_17_buffer[!clk]) ||(PRED7_18_buffer[clk] != PRED7_18_buffer[!clk]) ||(PRED7_19_buffer[clk] != PRED7_19_buffer[!clk]) ||(PRED7_20_buffer[clk] != PRED7_20_buffer[!clk]) ||(PRED7_21_buffer[clk] != PRED7_21_buffer[!clk]) ||(PRED7_22_buffer[clk] != PRED7_22_buffer[!clk]) ||(PRED7_23_buffer[clk] != PRED7_23_buffer[!clk]) ||(PRED7_24_buffer[clk] != PRED7_24_buffer[!clk]) ||(PRED7_25_buffer[clk] != PRED7_25_buffer[!clk]) ||(PRED7_26_buffer[clk] != PRED7_26_buffer[!clk]) ||(PRED7_27_buffer[clk] != PRED7_27_buffer[!clk]) ||(PRED7_28_buffer[clk] != PRED7_28_buffer[!clk]) ||(PRED7_29_buffer[clk] != PRED7_29_buffer[!clk]) ||(PRED7_30_buffer[clk] != PRED7_30_buffer[!clk]) ||(PRED7_31_buffer[clk] != PRED7_31_buffer[!clk]) ||(PRED15_0_buffer[clk] != PRED15_0_buffer[!clk]) ||(PRED15_1_buffer[clk] != PRED15_1_buffer[!clk]) ||(PRED15_2_buffer[clk] != PRED15_2_buffer[!clk]) ||(PRED15_3_buffer[clk] != PRED15_3_buffer[!clk]) ||(PRED15_4_buffer[clk] != PRED15_4_buffer[!clk]) ||(PRED15_5_buffer[clk] != PRED15_5_buffer[!clk]) ||(PRED15_6_buffer[clk] != PRED15_6_buffer[!clk]) ||(PRED15_7_buffer[clk] != PRED15_7_buffer[!clk]) ||(PRED15_8_buffer[clk] != PRED15_8_buffer[!clk]) ||(PRED15_9_buffer[clk] != PRED15_9_buffer[!clk]) ||(PRED15_10_buffer[clk] != PRED15_10_buffer[!clk]) ||(PRED15_11_buffer[clk] != PRED15_11_buffer[!clk]) ||(PRED15_12_buffer[clk] != PRED15_12_buffer[!clk]) ||(PRED15_13_buffer[clk] != PRED15_13_buffer[!clk]) ||(PRED15_14_buffer[clk] != PRED15_14_buffer[!clk]) ||(PRED15_15_buffer[clk] != PRED15_15_buffer[!clk]) ||(PRED15_16_buffer[clk] != PRED15_16_buffer[!clk]) ||(PRED15_17_buffer[clk] != PRED15_17_buffer[!clk]) ||(PRED15_18_buffer[clk] != PRED15_18_buffer[!clk]) ||(PRED15_19_buffer[clk] != PRED15_19_buffer[!clk]) ||(PRED15_20_buffer[clk] != PRED15_20_buffer[!clk]) ||(PRED15_21_buffer[clk] != PRED15_21_buffer[!clk]) ||(PRED15_22_buffer[clk] != PRED15_22_buffer[!clk]) ||(PRED15_23_buffer[clk] != PRED15_23_buffer[!clk]) ||(PRED15_24_buffer[clk] != PRED15_24_buffer[!clk]) ||(PRED15_25_buffer[clk] != PRED15_25_buffer[!clk]) ||(PRED15_26_buffer[clk] != PRED15_26_buffer[!clk]) ||(PRED15_27_buffer[clk] != PRED15_27_buffer[!clk]) ||(PRED15_28_buffer[clk] != PRED15_28_buffer[!clk]) ||(PRED15_29_buffer[clk] != PRED15_29_buffer[!clk]) ||(PRED15_30_buffer[clk] != PRED15_30_buffer[!clk]) ||(PRED15_31_buffer[clk] != PRED15_31_buffer[!clk]) ||(PRED23_0_buffer[clk] != PRED23_0_buffer[!clk]) ||(PRED23_1_buffer[clk] != PRED23_1_buffer[!clk]) ||(PRED23_2_buffer[clk] != PRED23_2_buffer[!clk]) ||(PRED23_3_buffer[clk] != PRED23_3_buffer[!clk]) ||(PRED23_4_buffer[clk] != PRED23_4_buffer[!clk]) ||(PRED23_5_buffer[clk] != PRED23_5_buffer[!clk]) ||(PRED23_6_buffer[clk] != PRED23_6_buffer[!clk]) ||(PRED23_7_buffer[clk] != PRED23_7_buffer[!clk]) ||(PRED23_8_buffer[clk] != PRED23_8_buffer[!clk]) ||(PRED23_9_buffer[clk] != PRED23_9_buffer[!clk]) ||(PRED23_10_buffer[clk] != PRED23_10_buffer[!clk]) ||(PRED23_11_buffer[clk] != PRED23_11_buffer[!clk]) ||(PRED23_12_buffer[clk] != PRED23_12_buffer[!clk]) ||(PRED23_13_buffer[clk] != PRED23_13_buffer[!clk]) ||(PRED23_14_buffer[clk] != PRED23_14_buffer[!clk]) ||(PRED23_15_buffer[clk] != PRED23_15_buffer[!clk]) ||(PRED23_16_buffer[clk] != PRED23_16_buffer[!clk]) ||(PRED23_17_buffer[clk] != PRED23_17_buffer[!clk]) ||(PRED23_18_buffer[clk] != PRED23_18_buffer[!clk]) ||(PRED23_19_buffer[clk] != PRED23_19_buffer[!clk]) ||(PRED23_20_buffer[clk] != PRED23_20_buffer[!clk]) ||(PRED23_21_buffer[clk] != PRED23_21_buffer[!clk]) ||(PRED23_22_buffer[clk] != PRED23_22_buffer[!clk]) ||(PRED23_23_buffer[clk] != PRED23_23_buffer[!clk]) ||(PRED23_24_buffer[clk] != PRED23_24_buffer[!clk]) ||(PRED23_25_buffer[clk] != PRED23_25_buffer[!clk]) ||(PRED23_26_buffer[clk] != PRED23_26_buffer[!clk]) ||(PRED23_27_buffer[clk] != PRED23_27_buffer[!clk]) ||(PRED23_28_buffer[clk] != PRED23_28_buffer[!clk]) ||(PRED23_29_buffer[clk] != PRED23_29_buffer[!clk]) ||(PRED23_30_buffer[clk] != PRED23_30_buffer[!clk]) ||(PRED23_31_buffer[clk] != PRED23_31_buffer[!clk]) ||(PRED31_0_buffer[clk] != PRED31_0_buffer[!clk]) ||(PRED31_1_buffer[clk] != PRED31_1_buffer[!clk]) ||(PRED31_2_buffer[clk] != PRED31_2_buffer[!clk]) ||(PRED31_3_buffer[clk] != PRED31_3_buffer[!clk]) ||(PRED31_4_buffer[clk] != PRED31_4_buffer[!clk]) ||(PRED31_5_buffer[clk] != PRED31_5_buffer[!clk]) ||(PRED31_6_buffer[clk] != PRED31_6_buffer[!clk]) ||(PRED31_7_buffer[clk] != PRED31_7_buffer[!clk]) ||(PRED31_8_buffer[clk] != PRED31_8_buffer[!clk]) ||(PRED31_9_buffer[clk] != PRED31_9_buffer[!clk]) ||(PRED31_10_buffer[clk] != PRED31_10_buffer[!clk]) ||(PRED31_11_buffer[clk] != PRED31_11_buffer[!clk]) ||(PRED31_12_buffer[clk] != PRED31_12_buffer[!clk]) ||(PRED31_13_buffer[clk] != PRED31_13_buffer[!clk]) ||(PRED31_14_buffer[clk] != PRED31_14_buffer[!clk]) ||(PRED31_15_buffer[clk] != PRED31_15_buffer[!clk]) ||(PRED31_16_buffer[clk] != PRED31_16_buffer[!clk]) ||(PRED31_17_buffer[clk] != PRED31_17_buffer[!clk]) ||(PRED31_18_buffer[clk] != PRED31_18_buffer[!clk]) ||(PRED31_19_buffer[clk] != PRED31_19_buffer[!clk]) ||(PRED31_20_buffer[clk] != PRED31_20_buffer[!clk]) ||(PRED31_21_buffer[clk] != PRED31_21_buffer[!clk]) ||(PRED31_22_buffer[clk] != PRED31_22_buffer[!clk]) ||(PRED31_23_buffer[clk] != PRED31_23_buffer[!clk]) ||(PRED31_24_buffer[clk] != PRED31_24_buffer[!clk]) ||(PRED31_25_buffer[clk] != PRED31_25_buffer[!clk]) ||(PRED31_26_buffer[clk] != PRED31_26_buffer[!clk]) ||(PRED31_27_buffer[clk] != PRED31_27_buffer[!clk]) ||(PRED31_28_buffer[clk] != PRED31_28_buffer[!clk]) ||(PRED31_29_buffer[clk] != PRED31_29_buffer[!clk]) ||(PRED31_30_buffer[clk] != PRED31_30_buffer[!clk]) ||(PRED31_31_buffer[clk] != PRED31_31_buffer[!clk]) ||(PRED39_0_buffer[clk] != PRED39_0_buffer[!clk]) ||(PRED39_1_buffer[clk] != PRED39_1_buffer[!clk]) ||(PRED39_2_buffer[clk] != PRED39_2_buffer[!clk]) ||(PRED39_3_buffer[clk] != PRED39_3_buffer[!clk]) ||(PRED39_4_buffer[clk] != PRED39_4_buffer[!clk]) ||(PRED39_5_buffer[clk] != PRED39_5_buffer[!clk]) ||(PRED39_6_buffer[clk] != PRED39_6_buffer[!clk]) ||(PRED39_7_buffer[clk] != PRED39_7_buffer[!clk]) ||(PRED39_8_buffer[clk] != PRED39_8_buffer[!clk]) ||(PRED39_9_buffer[clk] != PRED39_9_buffer[!clk]) ||(PRED39_10_buffer[clk] != PRED39_10_buffer[!clk]) ||(PRED39_11_buffer[clk] != PRED39_11_buffer[!clk]) ||(PRED39_12_buffer[clk] != PRED39_12_buffer[!clk]) ||(PRED39_13_buffer[clk] != PRED39_13_buffer[!clk]) ||(PRED39_14_buffer[clk] != PRED39_14_buffer[!clk]) ||(PRED39_15_buffer[clk] != PRED39_15_buffer[!clk]) ||(PRED39_16_buffer[clk] != PRED39_16_buffer[!clk]) ||(PRED39_17_buffer[clk] != PRED39_17_buffer[!clk]) ||(PRED39_18_buffer[clk] != PRED39_18_buffer[!clk]) ||(PRED39_19_buffer[clk] != PRED39_19_buffer[!clk]) ||(PRED39_20_buffer[clk] != PRED39_20_buffer[!clk]) ||(PRED39_21_buffer[clk] != PRED39_21_buffer[!clk]) ||(PRED39_22_buffer[clk] != PRED39_22_buffer[!clk]) ||(PRED39_23_buffer[clk] != PRED39_23_buffer[!clk]) ||(PRED39_24_buffer[clk] != PRED39_24_buffer[!clk]) ||(PRED39_25_buffer[clk] != PRED39_25_buffer[!clk]) ||(PRED39_26_buffer[clk] != PRED39_26_buffer[!clk]) ||(PRED39_27_buffer[clk] != PRED39_27_buffer[!clk]) ||(PRED39_28_buffer[clk] != PRED39_28_buffer[!clk]) ||(PRED39_29_buffer[clk] != PRED39_29_buffer[!clk]) ||(PRED39_30_buffer[clk] != PRED39_30_buffer[!clk]) ||(PRED39_31_buffer[clk] != PRED39_31_buffer[!clk]) ||(PRED47_0_buffer[clk] != PRED47_0_buffer[!clk]) ||(PRED47_1_buffer[clk] != PRED47_1_buffer[!clk]) ||(PRED47_2_buffer[clk] != PRED47_2_buffer[!clk]) ||(PRED47_3_buffer[clk] != PRED47_3_buffer[!clk]) ||(PRED47_4_buffer[clk] != PRED47_4_buffer[!clk]) ||(PRED47_5_buffer[clk] != PRED47_5_buffer[!clk]) ||(PRED47_6_buffer[clk] != PRED47_6_buffer[!clk]) ||(PRED47_7_buffer[clk] != PRED47_7_buffer[!clk]) ||(PRED47_8_buffer[clk] != PRED47_8_buffer[!clk]) ||(PRED47_9_buffer[clk] != PRED47_9_buffer[!clk]) ||(PRED47_10_buffer[clk] != PRED47_10_buffer[!clk]) ||(PRED47_11_buffer[clk] != PRED47_11_buffer[!clk]) ||(PRED47_12_buffer[clk] != PRED47_12_buffer[!clk]) ||(PRED47_13_buffer[clk] != PRED47_13_buffer[!clk]) ||(PRED47_14_buffer[clk] != PRED47_14_buffer[!clk]) ||(PRED47_15_buffer[clk] != PRED47_15_buffer[!clk]) ||(PRED47_16_buffer[clk] != PRED47_16_buffer[!clk]) ||(PRED47_17_buffer[clk] != PRED47_17_buffer[!clk]) ||(PRED47_18_buffer[clk] != PRED47_18_buffer[!clk]) ||(PRED47_19_buffer[clk] != PRED47_19_buffer[!clk]) ||(PRED47_20_buffer[clk] != PRED47_20_buffer[!clk]) ||(PRED47_21_buffer[clk] != PRED47_21_buffer[!clk]) ||(PRED47_22_buffer[clk] != PRED47_22_buffer[!clk]) ||(PRED47_23_buffer[clk] != PRED47_23_buffer[!clk]) ||(PRED47_24_buffer[clk] != PRED47_24_buffer[!clk]) ||(PRED47_25_buffer[clk] != PRED47_25_buffer[!clk]) ||(PRED47_26_buffer[clk] != PRED47_26_buffer[!clk]) ||(PRED47_27_buffer[clk] != PRED47_27_buffer[!clk]) ||(PRED47_28_buffer[clk] != PRED47_28_buffer[!clk]) ||(PRED47_29_buffer[clk] != PRED47_29_buffer[!clk]) ||(PRED47_30_buffer[clk] != PRED47_30_buffer[!clk]) ||(PRED47_31_buffer[clk] != PRED47_31_buffer[!clk]) ||(PRED55_0_buffer[clk] != PRED55_0_buffer[!clk]) ||(PRED55_1_buffer[clk] != PRED55_1_buffer[!clk]) ||(PRED55_2_buffer[clk] != PRED55_2_buffer[!clk]) ||(PRED55_3_buffer[clk] != PRED55_3_buffer[!clk]) ||(PRED55_4_buffer[clk] != PRED55_4_buffer[!clk]) ||(PRED55_5_buffer[clk] != PRED55_5_buffer[!clk]) ||(PRED55_6_buffer[clk] != PRED55_6_buffer[!clk]) ||(PRED55_7_buffer[clk] != PRED55_7_buffer[!clk]) ||(PRED55_8_buffer[clk] != PRED55_8_buffer[!clk]) ||(PRED55_9_buffer[clk] != PRED55_9_buffer[!clk]) ||(PRED55_10_buffer[clk] != PRED55_10_buffer[!clk]) ||(PRED55_11_buffer[clk] != PRED55_11_buffer[!clk]) ||(PRED55_12_buffer[clk] != PRED55_12_buffer[!clk]) ||(PRED55_13_buffer[clk] != PRED55_13_buffer[!clk]) ||(PRED55_14_buffer[clk] != PRED55_14_buffer[!clk]) ||(PRED55_15_buffer[clk] != PRED55_15_buffer[!clk]) ||(PRED55_16_buffer[clk] != PRED55_16_buffer[!clk]) ||(PRED55_17_buffer[clk] != PRED55_17_buffer[!clk]) ||(PRED55_18_buffer[clk] != PRED55_18_buffer[!clk]) ||(PRED55_19_buffer[clk] != PRED55_19_buffer[!clk]) ||(PRED55_20_buffer[clk] != PRED55_20_buffer[!clk]) ||(PRED55_21_buffer[clk] != PRED55_21_buffer[!clk]) ||(PRED55_22_buffer[clk] != PRED55_22_buffer[!clk]) ||(PRED55_23_buffer[clk] != PRED55_23_buffer[!clk]) ||(PRED55_24_buffer[clk] != PRED55_24_buffer[!clk]) ||(PRED55_25_buffer[clk] != PRED55_25_buffer[!clk]) ||(PRED55_26_buffer[clk] != PRED55_26_buffer[!clk]) ||(PRED55_27_buffer[clk] != PRED55_27_buffer[!clk]) ||(PRED55_28_buffer[clk] != PRED55_28_buffer[!clk]) ||(PRED55_29_buffer[clk] != PRED55_29_buffer[!clk]) ||(PRED55_30_buffer[clk] != PRED55_30_buffer[!clk]) ||(PRED55_31_buffer[clk] != PRED55_31_buffer[!clk]) ||(PRED63_0_buffer[clk] != PRED63_0_buffer[!clk]) ||(PRED63_1_buffer[clk] != PRED63_1_buffer[!clk]) ||(PRED63_2_buffer[clk] != PRED63_2_buffer[!clk]) ||(PRED63_3_buffer[clk] != PRED63_3_buffer[!clk]) ||(PRED63_4_buffer[clk] != PRED63_4_buffer[!clk]) ||(PRED63_5_buffer[clk] != PRED63_5_buffer[!clk]) ||(PRED63_6_buffer[clk] != PRED63_6_buffer[!clk]) ||(PRED63_7_buffer[clk] != PRED63_7_buffer[!clk]) ||(PRED63_8_buffer[clk] != PRED63_8_buffer[!clk]) ||(PRED63_9_buffer[clk] != PRED63_9_buffer[!clk]) ||(PRED63_10_buffer[clk] != PRED63_10_buffer[!clk]) ||(PRED63_11_buffer[clk] != PRED63_11_buffer[!clk]) ||(PRED63_12_buffer[clk] != PRED63_12_buffer[!clk]) ||(PRED63_13_buffer[clk] != PRED63_13_buffer[!clk]) ||(PRED63_14_buffer[clk] != PRED63_14_buffer[!clk]) ||(PRED63_15_buffer[clk] != PRED63_15_buffer[!clk]) ||(PRED63_16_buffer[clk] != PRED63_16_buffer[!clk]) ||(PRED63_17_buffer[clk] != PRED63_17_buffer[!clk]) ||(PRED63_18_buffer[clk] != PRED63_18_buffer[!clk]) ||(PRED63_19_buffer[clk] != PRED63_19_buffer[!clk]) ||(PRED63_20_buffer[clk] != PRED63_20_buffer[!clk]) ||(PRED63_21_buffer[clk] != PRED63_21_buffer[!clk]) ||(PRED63_22_buffer[clk] != PRED63_22_buffer[!clk]) ||(PRED63_23_buffer[clk] != PRED63_23_buffer[!clk]) ||(PRED63_24_buffer[clk] != PRED63_24_buffer[!clk]) ||(PRED63_25_buffer[clk] != PRED63_25_buffer[!clk]) ||(PRED63_26_buffer[clk] != PRED63_26_buffer[!clk]) ||(PRED63_27_buffer[clk] != PRED63_27_buffer[!clk]) ||(PRED63_28_buffer[clk] != PRED63_28_buffer[!clk]) ||(PRED63_29_buffer[clk] != PRED63_29_buffer[!clk]) ||(PRED63_30_buffer[clk] != PRED63_30_buffer[!clk]) ||(PRED63_31_buffer[clk] != PRED63_31_buffer[!clk]) ) begin
      warp7_sig = 1'b1;
    end else begin
      warp7_sig = 1'b0;
    end

  end

  // Determine if there is a change in any of the register files
  // When there is a change, then print out the statements below

  // Need to add timestamp, PC start, PC finish, all of Warp Data
  // Output Register Changes
  initial begin
    for (i = 0 ; i < 10000 ; i = i + 1) begin
      @ (posedge clk);
      // pick which warp to trace // WARPEDIT
      if ( warp7_sig == 1'b1 ) begin // change warpX_sig to select
        $fwrite(f, " \n=====================================================\n");
        $fwrite(f, "Simulation Time          ---> ", $time);
        $fwrite(f, "\n\n");

        if (PRED0_0_buffer[clk] != PRED0_0_buffer[!clk]) begin
          $fwrite(f, "Register (0,0) Value: %h\n", PRED0_0_buffer[clk]);
        end
        if (PRED0_1_buffer[clk] != PRED0_1_buffer[!clk]) begin
          $fwrite(f, "Register (0,1) Value: %h\n", PRED0_1_buffer[clk]);
        end
        if (PRED0_2_buffer[clk] != PRED0_2_buffer[!clk]) begin
          $fwrite(f, "Register (0,2) Value: %h\n", PRED0_2_buffer[clk]);
        end
        if (PRED0_3_buffer[clk] != PRED0_3_buffer[!clk]) begin
          $fwrite(f, "Register (0,3) Value: %h\n", PRED0_3_buffer[clk]);
        end
        if (PRED0_4_buffer[clk] != PRED0_4_buffer[!clk]) begin
          $fwrite(f, "Register (0,4) Value: %h\n", PRED0_4_buffer[clk]);
        end
        if (PRED0_5_buffer[clk] != PRED0_5_buffer[!clk]) begin
          $fwrite(f, "Register (0,5) Value: %h\n", PRED0_5_buffer[clk]);
        end
        if (PRED0_6_buffer[clk] != PRED0_6_buffer[!clk]) begin
          $fwrite(f, "Register (0,6) Value: %h\n", PRED0_6_buffer[clk]);
        end
        if (PRED0_7_buffer[clk] != PRED0_7_buffer[!clk]) begin
          $fwrite(f, "Register (0,7) Value: %h\n", PRED0_7_buffer[clk]);
        end
        if (PRED0_8_buffer[clk] != PRED0_8_buffer[!clk]) begin
          $fwrite(f, "Register (0,8) Value: %h\n", PRED0_8_buffer[clk]);
        end
        if (PRED0_9_buffer[clk] != PRED0_9_buffer[!clk]) begin
          $fwrite(f, "Register (0,9) Value: %h\n", PRED0_9_buffer[clk]);
        end
        if (PRED0_10_buffer[clk] != PRED0_10_buffer[!clk]) begin
          $fwrite(f, "Register (0,10) Value: %h\n", PRED0_10_buffer[clk]);
        end
        if (PRED0_11_buffer[clk] != PRED0_11_buffer[!clk]) begin
          $fwrite(f, "Register (0,11) Value: %h\n", PRED0_11_buffer[clk]);
        end
        if (PRED0_12_buffer[clk] != PRED0_12_buffer[!clk]) begin
          $fwrite(f, "Register (0,12) Value: %h\n", PRED0_12_buffer[clk]);
        end
        if (PRED0_13_buffer[clk] != PRED0_13_buffer[!clk]) begin
          $fwrite(f, "Register (0,13) Value: %h\n", PRED0_13_buffer[clk]);
        end
        if (PRED0_14_buffer[clk] != PRED0_14_buffer[!clk]) begin
          $fwrite(f, "Register (0,14) Value: %h\n", PRED0_14_buffer[clk]);
        end
        if (PRED0_15_buffer[clk] != PRED0_15_buffer[!clk]) begin
          $fwrite(f, "Register (0,15) Value: %h\n", PRED0_15_buffer[clk]);
        end
        if (PRED0_16_buffer[clk] != PRED0_16_buffer[!clk]) begin
          $fwrite(f, "Register (0,16) Value: %h\n", PRED0_16_buffer[clk]);
        end
        if (PRED0_17_buffer[clk] != PRED0_17_buffer[!clk]) begin
          $fwrite(f, "Register (0,17) Value: %h\n", PRED0_17_buffer[clk]);
        end
        if (PRED0_18_buffer[clk] != PRED0_18_buffer[!clk]) begin
          $fwrite(f, "Register (0,18) Value: %h\n", PRED0_18_buffer[clk]);
        end
        if (PRED0_19_buffer[clk] != PRED0_19_buffer[!clk]) begin
          $fwrite(f, "Register (0,19) Value: %h\n", PRED0_19_buffer[clk]);
        end
        if (PRED0_20_buffer[clk] != PRED0_20_buffer[!clk]) begin
          $fwrite(f, "Register (0,20) Value: %h\n", PRED0_20_buffer[clk]);
        end
        if (PRED0_21_buffer[clk] != PRED0_21_buffer[!clk]) begin
          $fwrite(f, "Register (0,21) Value: %h\n", PRED0_21_buffer[clk]);
        end
        if (PRED0_22_buffer[clk] != PRED0_22_buffer[!clk]) begin
          $fwrite(f, "Register (0,22) Value: %h\n", PRED0_22_buffer[clk]);
        end
        if (PRED0_23_buffer[clk] != PRED0_23_buffer[!clk]) begin
          $fwrite(f, "Register (0,23) Value: %h\n", PRED0_23_buffer[clk]);
        end
        if (PRED0_24_buffer[clk] != PRED0_24_buffer[!clk]) begin
          $fwrite(f, "Register (0,24) Value: %h\n", PRED0_24_buffer[clk]);
        end
        if (PRED0_25_buffer[clk] != PRED0_25_buffer[!clk]) begin
          $fwrite(f, "Register (0,25) Value: %h\n", PRED0_25_buffer[clk]);
        end
        if (PRED0_26_buffer[clk] != PRED0_26_buffer[!clk]) begin
          $fwrite(f, "Register (0,26) Value: %h\n", PRED0_26_buffer[clk]);
        end
        if (PRED0_27_buffer[clk] != PRED0_27_buffer[!clk]) begin
          $fwrite(f, "Register (0,27) Value: %h\n", PRED0_27_buffer[clk]);
        end
        if (PRED0_28_buffer[clk] != PRED0_28_buffer[!clk]) begin
          $fwrite(f, "Register (0,28) Value: %h\n", PRED0_28_buffer[clk]);
        end
        if (PRED0_29_buffer[clk] != PRED0_29_buffer[!clk]) begin
          $fwrite(f, "Register (0,29) Value: %h\n", PRED0_29_buffer[clk]);
        end
        if (PRED0_30_buffer[clk] != PRED0_30_buffer[!clk]) begin
          $fwrite(f, "Register (0,30) Value: %h\n", PRED0_30_buffer[clk]);
        end
        if (PRED0_31_buffer[clk] != PRED0_31_buffer[!clk]) begin
          $fwrite(f, "Register (0,31) Value: %h\n", PRED0_31_buffer[clk]);
        end
        if (PRED1_0_buffer[clk] != PRED1_0_buffer[!clk]) begin
          $fwrite(f, "Register (1,0) Value: %h\n", PRED1_0_buffer[clk]);
        end
        if (PRED1_1_buffer[clk] != PRED1_1_buffer[!clk]) begin
          $fwrite(f, "Register (1,1) Value: %h\n", PRED1_1_buffer[clk]);
        end
        if (PRED1_2_buffer[clk] != PRED1_2_buffer[!clk]) begin
          $fwrite(f, "Register (1,2) Value: %h\n", PRED1_2_buffer[clk]);
        end
        if (PRED1_3_buffer[clk] != PRED1_3_buffer[!clk]) begin
          $fwrite(f, "Register (1,3) Value: %h\n", PRED1_3_buffer[clk]);
        end
        if (PRED1_4_buffer[clk] != PRED1_4_buffer[!clk]) begin
          $fwrite(f, "Register (1,4) Value: %h\n", PRED1_4_buffer[clk]);
        end
        if (PRED1_5_buffer[clk] != PRED1_5_buffer[!clk]) begin
          $fwrite(f, "Register (1,5) Value: %h\n", PRED1_5_buffer[clk]);
        end
        if (PRED1_6_buffer[clk] != PRED1_6_buffer[!clk]) begin
          $fwrite(f, "Register (1,6) Value: %h\n", PRED1_6_buffer[clk]);
        end
        if (PRED1_7_buffer[clk] != PRED1_7_buffer[!clk]) begin
          $fwrite(f, "Register (1,7) Value: %h\n", PRED1_7_buffer[clk]);
        end
        if (PRED1_8_buffer[clk] != PRED1_8_buffer[!clk]) begin
          $fwrite(f, "Register (1,8) Value: %h\n", PRED1_8_buffer[clk]);
        end
        if (PRED1_9_buffer[clk] != PRED1_9_buffer[!clk]) begin
          $fwrite(f, "Register (1,9) Value: %h\n", PRED1_9_buffer[clk]);
        end
        if (PRED1_10_buffer[clk] != PRED1_10_buffer[!clk]) begin
          $fwrite(f, "Register (1,10) Value: %h\n", PRED1_10_buffer[clk]);
        end
        if (PRED1_11_buffer[clk] != PRED1_11_buffer[!clk]) begin
          $fwrite(f, "Register (1,11) Value: %h\n", PRED1_11_buffer[clk]);
        end
        if (PRED1_12_buffer[clk] != PRED1_12_buffer[!clk]) begin
          $fwrite(f, "Register (1,12) Value: %h\n", PRED1_12_buffer[clk]);
        end
        if (PRED1_13_buffer[clk] != PRED1_13_buffer[!clk]) begin
          $fwrite(f, "Register (1,13) Value: %h\n", PRED1_13_buffer[clk]);
        end
        if (PRED1_14_buffer[clk] != PRED1_14_buffer[!clk]) begin
          $fwrite(f, "Register (1,14) Value: %h\n", PRED1_14_buffer[clk]);
        end
        if (PRED1_15_buffer[clk] != PRED1_15_buffer[!clk]) begin
          $fwrite(f, "Register (1,15) Value: %h\n", PRED1_15_buffer[clk]);
        end
        if (PRED1_16_buffer[clk] != PRED1_16_buffer[!clk]) begin
          $fwrite(f, "Register (1,16) Value: %h\n", PRED1_16_buffer[clk]);
        end
        if (PRED1_17_buffer[clk] != PRED1_17_buffer[!clk]) begin
          $fwrite(f, "Register (1,17) Value: %h\n", PRED1_17_buffer[clk]);
        end
        if (PRED1_18_buffer[clk] != PRED1_18_buffer[!clk]) begin
          $fwrite(f, "Register (1,18) Value: %h\n", PRED1_18_buffer[clk]);
        end
        if (PRED1_19_buffer[clk] != PRED1_19_buffer[!clk]) begin
          $fwrite(f, "Register (1,19) Value: %h\n", PRED1_19_buffer[clk]);
        end
        if (PRED1_20_buffer[clk] != PRED1_20_buffer[!clk]) begin
          $fwrite(f, "Register (1,20) Value: %h\n", PRED1_20_buffer[clk]);
        end
        if (PRED1_21_buffer[clk] != PRED1_21_buffer[!clk]) begin
          $fwrite(f, "Register (1,21) Value: %h\n", PRED1_21_buffer[clk]);
        end
        if (PRED1_22_buffer[clk] != PRED1_22_buffer[!clk]) begin
          $fwrite(f, "Register (1,22) Value: %h\n", PRED1_22_buffer[clk]);
        end
        if (PRED1_23_buffer[clk] != PRED1_23_buffer[!clk]) begin
          $fwrite(f, "Register (1,23) Value: %h\n", PRED1_23_buffer[clk]);
        end
        if (PRED1_24_buffer[clk] != PRED1_24_buffer[!clk]) begin
          $fwrite(f, "Register (1,24) Value: %h\n", PRED1_24_buffer[clk]);
        end
        if (PRED1_25_buffer[clk] != PRED1_25_buffer[!clk]) begin
          $fwrite(f, "Register (1,25) Value: %h\n", PRED1_25_buffer[clk]);
        end
        if (PRED1_26_buffer[clk] != PRED1_26_buffer[!clk]) begin
          $fwrite(f, "Register (1,26) Value: %h\n", PRED1_26_buffer[clk]);
        end
        if (PRED1_27_buffer[clk] != PRED1_27_buffer[!clk]) begin
          $fwrite(f, "Register (1,27) Value: %h\n", PRED1_27_buffer[clk]);
        end
        if (PRED1_28_buffer[clk] != PRED1_28_buffer[!clk]) begin
          $fwrite(f, "Register (1,28) Value: %h\n", PRED1_28_buffer[clk]);
        end
        if (PRED1_29_buffer[clk] != PRED1_29_buffer[!clk]) begin
          $fwrite(f, "Register (1,29) Value: %h\n", PRED1_29_buffer[clk]);
        end
        if (PRED1_30_buffer[clk] != PRED1_30_buffer[!clk]) begin
          $fwrite(f, "Register (1,30) Value: %h\n", PRED1_30_buffer[clk]);
        end
        if (PRED1_31_buffer[clk] != PRED1_31_buffer[!clk]) begin
          $fwrite(f, "Register (1,31) Value: %h\n", PRED1_31_buffer[clk]);
        end
        if (PRED2_0_buffer[clk] != PRED2_0_buffer[!clk]) begin
          $fwrite(f, "Register (2,0) Value: %h\n", PRED2_0_buffer[clk]);
        end
        if (PRED2_1_buffer[clk] != PRED2_1_buffer[!clk]) begin
          $fwrite(f, "Register (2,1) Value: %h\n", PRED2_1_buffer[clk]);
        end
        if (PRED2_2_buffer[clk] != PRED2_2_buffer[!clk]) begin
          $fwrite(f, "Register (2,2) Value: %h\n", PRED2_2_buffer[clk]);
        end
        if (PRED2_3_buffer[clk] != PRED2_3_buffer[!clk]) begin
          $fwrite(f, "Register (2,3) Value: %h\n", PRED2_3_buffer[clk]);
        end
        if (PRED2_4_buffer[clk] != PRED2_4_buffer[!clk]) begin
          $fwrite(f, "Register (2,4) Value: %h\n", PRED2_4_buffer[clk]);
        end
        if (PRED2_5_buffer[clk] != PRED2_5_buffer[!clk]) begin
          $fwrite(f, "Register (2,5) Value: %h\n", PRED2_5_buffer[clk]);
        end
        if (PRED2_6_buffer[clk] != PRED2_6_buffer[!clk]) begin
          $fwrite(f, "Register (2,6) Value: %h\n", PRED2_6_buffer[clk]);
        end
        if (PRED2_7_buffer[clk] != PRED2_7_buffer[!clk]) begin
          $fwrite(f, "Register (2,7) Value: %h\n", PRED2_7_buffer[clk]);
        end
        if (PRED2_8_buffer[clk] != PRED2_8_buffer[!clk]) begin
          $fwrite(f, "Register (2,8) Value: %h\n", PRED2_8_buffer[clk]);
        end
        if (PRED2_9_buffer[clk] != PRED2_9_buffer[!clk]) begin
          $fwrite(f, "Register (2,9) Value: %h\n", PRED2_9_buffer[clk]);
        end
        if (PRED2_10_buffer[clk] != PRED2_10_buffer[!clk]) begin
          $fwrite(f, "Register (2,10) Value: %h\n", PRED2_10_buffer[clk]);
        end
        if (PRED2_11_buffer[clk] != PRED2_11_buffer[!clk]) begin
          $fwrite(f, "Register (2,11) Value: %h\n", PRED2_11_buffer[clk]);
        end
        if (PRED2_12_buffer[clk] != PRED2_12_buffer[!clk]) begin
          $fwrite(f, "Register (2,12) Value: %h\n", PRED2_12_buffer[clk]);
        end
        if (PRED2_13_buffer[clk] != PRED2_13_buffer[!clk]) begin
          $fwrite(f, "Register (2,13) Value: %h\n", PRED2_13_buffer[clk]);
        end
        if (PRED2_14_buffer[clk] != PRED2_14_buffer[!clk]) begin
          $fwrite(f, "Register (2,14) Value: %h\n", PRED2_14_buffer[clk]);
        end
        if (PRED2_15_buffer[clk] != PRED2_15_buffer[!clk]) begin
          $fwrite(f, "Register (2,15) Value: %h\n", PRED2_15_buffer[clk]);
        end
        if (PRED2_16_buffer[clk] != PRED2_16_buffer[!clk]) begin
          $fwrite(f, "Register (2,16) Value: %h\n", PRED2_16_buffer[clk]);
        end
        if (PRED2_17_buffer[clk] != PRED2_17_buffer[!clk]) begin
          $fwrite(f, "Register (2,17) Value: %h\n", PRED2_17_buffer[clk]);
        end
        if (PRED2_18_buffer[clk] != PRED2_18_buffer[!clk]) begin
          $fwrite(f, "Register (2,18) Value: %h\n", PRED2_18_buffer[clk]);
        end
        if (PRED2_19_buffer[clk] != PRED2_19_buffer[!clk]) begin
          $fwrite(f, "Register (2,19) Value: %h\n", PRED2_19_buffer[clk]);
        end
        if (PRED2_20_buffer[clk] != PRED2_20_buffer[!clk]) begin
          $fwrite(f, "Register (2,20) Value: %h\n", PRED2_20_buffer[clk]);
        end
        if (PRED2_21_buffer[clk] != PRED2_21_buffer[!clk]) begin
          $fwrite(f, "Register (2,21) Value: %h\n", PRED2_21_buffer[clk]);
        end
        if (PRED2_22_buffer[clk] != PRED2_22_buffer[!clk]) begin
          $fwrite(f, "Register (2,22) Value: %h\n", PRED2_22_buffer[clk]);
        end
        if (PRED2_23_buffer[clk] != PRED2_23_buffer[!clk]) begin
          $fwrite(f, "Register (2,23) Value: %h\n", PRED2_23_buffer[clk]);
        end
        if (PRED2_24_buffer[clk] != PRED2_24_buffer[!clk]) begin
          $fwrite(f, "Register (2,24) Value: %h\n", PRED2_24_buffer[clk]);
        end
        if (PRED2_25_buffer[clk] != PRED2_25_buffer[!clk]) begin
          $fwrite(f, "Register (2,25) Value: %h\n", PRED2_25_buffer[clk]);
        end
        if (PRED2_26_buffer[clk] != PRED2_26_buffer[!clk]) begin
          $fwrite(f, "Register (2,26) Value: %h\n", PRED2_26_buffer[clk]);
        end
        if (PRED2_27_buffer[clk] != PRED2_27_buffer[!clk]) begin
          $fwrite(f, "Register (2,27) Value: %h\n", PRED2_27_buffer[clk]);
        end
        if (PRED2_28_buffer[clk] != PRED2_28_buffer[!clk]) begin
          $fwrite(f, "Register (2,28) Value: %h\n", PRED2_28_buffer[clk]);
        end
        if (PRED2_29_buffer[clk] != PRED2_29_buffer[!clk]) begin
          $fwrite(f, "Register (2,29) Value: %h\n", PRED2_29_buffer[clk]);
        end
        if (PRED2_30_buffer[clk] != PRED2_30_buffer[!clk]) begin
          $fwrite(f, "Register (2,30) Value: %h\n", PRED2_30_buffer[clk]);
        end
        if (PRED2_31_buffer[clk] != PRED2_31_buffer[!clk]) begin
          $fwrite(f, "Register (2,31) Value: %h\n", PRED2_31_buffer[clk]);
        end
        if (PRED3_0_buffer[clk] != PRED3_0_buffer[!clk]) begin
          $fwrite(f, "Register (3,0) Value: %h\n", PRED3_0_buffer[clk]);
        end
        if (PRED3_1_buffer[clk] != PRED3_1_buffer[!clk]) begin
          $fwrite(f, "Register (3,1) Value: %h\n", PRED3_1_buffer[clk]);
        end
        if (PRED3_2_buffer[clk] != PRED3_2_buffer[!clk]) begin
          $fwrite(f, "Register (3,2) Value: %h\n", PRED3_2_buffer[clk]);
        end
        if (PRED3_3_buffer[clk] != PRED3_3_buffer[!clk]) begin
          $fwrite(f, "Register (3,3) Value: %h\n", PRED3_3_buffer[clk]);
        end
        if (PRED3_4_buffer[clk] != PRED3_4_buffer[!clk]) begin
          $fwrite(f, "Register (3,4) Value: %h\n", PRED3_4_buffer[clk]);
        end
        if (PRED3_5_buffer[clk] != PRED3_5_buffer[!clk]) begin
          $fwrite(f, "Register (3,5) Value: %h\n", PRED3_5_buffer[clk]);
        end
        if (PRED3_6_buffer[clk] != PRED3_6_buffer[!clk]) begin
          $fwrite(f, "Register (3,6) Value: %h\n", PRED3_6_buffer[clk]);
        end
        if (PRED3_7_buffer[clk] != PRED3_7_buffer[!clk]) begin
          $fwrite(f, "Register (3,7) Value: %h\n", PRED3_7_buffer[clk]);
        end
        if (PRED3_8_buffer[clk] != PRED3_8_buffer[!clk]) begin
          $fwrite(f, "Register (3,8) Value: %h\n", PRED3_8_buffer[clk]);
        end
        if (PRED3_9_buffer[clk] != PRED3_9_buffer[!clk]) begin
          $fwrite(f, "Register (3,9) Value: %h\n", PRED3_9_buffer[clk]);
        end
        if (PRED3_10_buffer[clk] != PRED3_10_buffer[!clk]) begin
          $fwrite(f, "Register (3,10) Value: %h\n", PRED3_10_buffer[clk]);
        end
        if (PRED3_11_buffer[clk] != PRED3_11_buffer[!clk]) begin
          $fwrite(f, "Register (3,11) Value: %h\n", PRED3_11_buffer[clk]);
        end
        if (PRED3_12_buffer[clk] != PRED3_12_buffer[!clk]) begin
          $fwrite(f, "Register (3,12) Value: %h\n", PRED3_12_buffer[clk]);
        end
        if (PRED3_13_buffer[clk] != PRED3_13_buffer[!clk]) begin
          $fwrite(f, "Register (3,13) Value: %h\n", PRED3_13_buffer[clk]);
        end
        if (PRED3_14_buffer[clk] != PRED3_14_buffer[!clk]) begin
          $fwrite(f, "Register (3,14) Value: %h\n", PRED3_14_buffer[clk]);
        end
        if (PRED3_15_buffer[clk] != PRED3_15_buffer[!clk]) begin
          $fwrite(f, "Register (3,15) Value: %h\n", PRED3_15_buffer[clk]);
        end
        if (PRED3_16_buffer[clk] != PRED3_16_buffer[!clk]) begin
          $fwrite(f, "Register (3,16) Value: %h\n", PRED3_16_buffer[clk]);
        end
        if (PRED3_17_buffer[clk] != PRED3_17_buffer[!clk]) begin
          $fwrite(f, "Register (3,17) Value: %h\n", PRED3_17_buffer[clk]);
        end
        if (PRED3_18_buffer[clk] != PRED3_18_buffer[!clk]) begin
          $fwrite(f, "Register (3,18) Value: %h\n", PRED3_18_buffer[clk]);
        end
        if (PRED3_19_buffer[clk] != PRED3_19_buffer[!clk]) begin
          $fwrite(f, "Register (3,19) Value: %h\n", PRED3_19_buffer[clk]);
        end
        if (PRED3_20_buffer[clk] != PRED3_20_buffer[!clk]) begin
          $fwrite(f, "Register (3,20) Value: %h\n", PRED3_20_buffer[clk]);
        end
        if (PRED3_21_buffer[clk] != PRED3_21_buffer[!clk]) begin
          $fwrite(f, "Register (3,21) Value: %h\n", PRED3_21_buffer[clk]);
        end
        if (PRED3_22_buffer[clk] != PRED3_22_buffer[!clk]) begin
          $fwrite(f, "Register (3,22) Value: %h\n", PRED3_22_buffer[clk]);
        end
        if (PRED3_23_buffer[clk] != PRED3_23_buffer[!clk]) begin
          $fwrite(f, "Register (3,23) Value: %h\n", PRED3_23_buffer[clk]);
        end
        if (PRED3_24_buffer[clk] != PRED3_24_buffer[!clk]) begin
          $fwrite(f, "Register (3,24) Value: %h\n", PRED3_24_buffer[clk]);
        end
        if (PRED3_25_buffer[clk] != PRED3_25_buffer[!clk]) begin
          $fwrite(f, "Register (3,25) Value: %h\n", PRED3_25_buffer[clk]);
        end
        if (PRED3_26_buffer[clk] != PRED3_26_buffer[!clk]) begin
          $fwrite(f, "Register (3,26) Value: %h\n", PRED3_26_buffer[clk]);
        end
        if (PRED3_27_buffer[clk] != PRED3_27_buffer[!clk]) begin
          $fwrite(f, "Register (3,27) Value: %h\n", PRED3_27_buffer[clk]);
        end
        if (PRED3_28_buffer[clk] != PRED3_28_buffer[!clk]) begin
          $fwrite(f, "Register (3,28) Value: %h\n", PRED3_28_buffer[clk]);
        end
        if (PRED3_29_buffer[clk] != PRED3_29_buffer[!clk]) begin
          $fwrite(f, "Register (3,29) Value: %h\n", PRED3_29_buffer[clk]);
        end
        if (PRED3_30_buffer[clk] != PRED3_30_buffer[!clk]) begin
          $fwrite(f, "Register (3,30) Value: %h\n", PRED3_30_buffer[clk]);
        end
        if (PRED3_31_buffer[clk] != PRED3_31_buffer[!clk]) begin
          $fwrite(f, "Register (3,31) Value: %h\n", PRED3_31_buffer[clk]);
        end
        if (PRED4_0_buffer[clk] != PRED4_0_buffer[!clk]) begin
          $fwrite(f, "Register (4,0) Value: %h\n", PRED4_0_buffer[clk]);
        end
        if (PRED4_1_buffer[clk] != PRED4_1_buffer[!clk]) begin
          $fwrite(f, "Register (4,1) Value: %h\n", PRED4_1_buffer[clk]);
        end
        if (PRED4_2_buffer[clk] != PRED4_2_buffer[!clk]) begin
          $fwrite(f, "Register (4,2) Value: %h\n", PRED4_2_buffer[clk]);
        end
        if (PRED4_3_buffer[clk] != PRED4_3_buffer[!clk]) begin
          $fwrite(f, "Register (4,3) Value: %h\n", PRED4_3_buffer[clk]);
        end
        if (PRED4_4_buffer[clk] != PRED4_4_buffer[!clk]) begin
          $fwrite(f, "Register (4,4) Value: %h\n", PRED4_4_buffer[clk]);
        end
        if (PRED4_5_buffer[clk] != PRED4_5_buffer[!clk]) begin
          $fwrite(f, "Register (4,5) Value: %h\n", PRED4_5_buffer[clk]);
        end
        if (PRED4_6_buffer[clk] != PRED4_6_buffer[!clk]) begin
          $fwrite(f, "Register (4,6) Value: %h\n", PRED4_6_buffer[clk]);
        end
        if (PRED4_7_buffer[clk] != PRED4_7_buffer[!clk]) begin
          $fwrite(f, "Register (4,7) Value: %h\n", PRED4_7_buffer[clk]);
        end
        if (PRED4_8_buffer[clk] != PRED4_8_buffer[!clk]) begin
          $fwrite(f, "Register (4,8) Value: %h\n", PRED4_8_buffer[clk]);
        end
        if (PRED4_9_buffer[clk] != PRED4_9_buffer[!clk]) begin
          $fwrite(f, "Register (4,9) Value: %h\n", PRED4_9_buffer[clk]);
        end
        if (PRED4_10_buffer[clk] != PRED4_10_buffer[!clk]) begin
          $fwrite(f, "Register (4,10) Value: %h\n", PRED4_10_buffer[clk]);
        end
        if (PRED4_11_buffer[clk] != PRED4_11_buffer[!clk]) begin
          $fwrite(f, "Register (4,11) Value: %h\n", PRED4_11_buffer[clk]);
        end
        if (PRED4_12_buffer[clk] != PRED4_12_buffer[!clk]) begin
          $fwrite(f, "Register (4,12) Value: %h\n", PRED4_12_buffer[clk]);
        end
        if (PRED4_13_buffer[clk] != PRED4_13_buffer[!clk]) begin
          $fwrite(f, "Register (4,13) Value: %h\n", PRED4_13_buffer[clk]);
        end
        if (PRED4_14_buffer[clk] != PRED4_14_buffer[!clk]) begin
          $fwrite(f, "Register (4,14) Value: %h\n", PRED4_14_buffer[clk]);
        end
        if (PRED4_15_buffer[clk] != PRED4_15_buffer[!clk]) begin
          $fwrite(f, "Register (4,15) Value: %h\n", PRED4_15_buffer[clk]);
        end
        if (PRED4_16_buffer[clk] != PRED4_16_buffer[!clk]) begin
          $fwrite(f, "Register (4,16) Value: %h\n", PRED4_16_buffer[clk]);
        end
        if (PRED4_17_buffer[clk] != PRED4_17_buffer[!clk]) begin
          $fwrite(f, "Register (4,17) Value: %h\n", PRED4_17_buffer[clk]);
        end
        if (PRED4_18_buffer[clk] != PRED4_18_buffer[!clk]) begin
          $fwrite(f, "Register (4,18) Value: %h\n", PRED4_18_buffer[clk]);
        end
        if (PRED4_19_buffer[clk] != PRED4_19_buffer[!clk]) begin
          $fwrite(f, "Register (4,19) Value: %h\n", PRED4_19_buffer[clk]);
        end
        if (PRED4_20_buffer[clk] != PRED4_20_buffer[!clk]) begin
          $fwrite(f, "Register (4,20) Value: %h\n", PRED4_20_buffer[clk]);
        end
        if (PRED4_21_buffer[clk] != PRED4_21_buffer[!clk]) begin
          $fwrite(f, "Register (4,21) Value: %h\n", PRED4_21_buffer[clk]);
        end
        if (PRED4_22_buffer[clk] != PRED4_22_buffer[!clk]) begin
          $fwrite(f, "Register (4,22) Value: %h\n", PRED4_22_buffer[clk]);
        end
        if (PRED4_23_buffer[clk] != PRED4_23_buffer[!clk]) begin
          $fwrite(f, "Register (4,23) Value: %h\n", PRED4_23_buffer[clk]);
        end
        if (PRED4_24_buffer[clk] != PRED4_24_buffer[!clk]) begin
          $fwrite(f, "Register (4,24) Value: %h\n", PRED4_24_buffer[clk]);
        end
        if (PRED4_25_buffer[clk] != PRED4_25_buffer[!clk]) begin
          $fwrite(f, "Register (4,25) Value: %h\n", PRED4_25_buffer[clk]);
        end
        if (PRED4_26_buffer[clk] != PRED4_26_buffer[!clk]) begin
          $fwrite(f, "Register (4,26) Value: %h\n", PRED4_26_buffer[clk]);
        end
        if (PRED4_27_buffer[clk] != PRED4_27_buffer[!clk]) begin
          $fwrite(f, "Register (4,27) Value: %h\n", PRED4_27_buffer[clk]);
        end
        if (PRED4_28_buffer[clk] != PRED4_28_buffer[!clk]) begin
          $fwrite(f, "Register (4,28) Value: %h\n", PRED4_28_buffer[clk]);
        end
        if (PRED4_29_buffer[clk] != PRED4_29_buffer[!clk]) begin
          $fwrite(f, "Register (4,29) Value: %h\n", PRED4_29_buffer[clk]);
        end
        if (PRED4_30_buffer[clk] != PRED4_30_buffer[!clk]) begin
          $fwrite(f, "Register (4,30) Value: %h\n", PRED4_30_buffer[clk]);
        end
        if (PRED4_31_buffer[clk] != PRED4_31_buffer[!clk]) begin
          $fwrite(f, "Register (4,31) Value: %h\n", PRED4_31_buffer[clk]);
        end
        if (PRED5_0_buffer[clk] != PRED5_0_buffer[!clk]) begin
          $fwrite(f, "Register (5,0) Value: %h\n", PRED5_0_buffer[clk]);
        end
        if (PRED5_1_buffer[clk] != PRED5_1_buffer[!clk]) begin
          $fwrite(f, "Register (5,1) Value: %h\n", PRED5_1_buffer[clk]);
        end
        if (PRED5_2_buffer[clk] != PRED5_2_buffer[!clk]) begin
          $fwrite(f, "Register (5,2) Value: %h\n", PRED5_2_buffer[clk]);
        end
        if (PRED5_3_buffer[clk] != PRED5_3_buffer[!clk]) begin
          $fwrite(f, "Register (5,3) Value: %h\n", PRED5_3_buffer[clk]);
        end
        if (PRED5_4_buffer[clk] != PRED5_4_buffer[!clk]) begin
          $fwrite(f, "Register (5,4) Value: %h\n", PRED5_4_buffer[clk]);
        end
        if (PRED5_5_buffer[clk] != PRED5_5_buffer[!clk]) begin
          $fwrite(f, "Register (5,5) Value: %h\n", PRED5_5_buffer[clk]);
        end
        if (PRED5_6_buffer[clk] != PRED5_6_buffer[!clk]) begin
          $fwrite(f, "Register (5,6) Value: %h\n", PRED5_6_buffer[clk]);
        end
        if (PRED5_7_buffer[clk] != PRED5_7_buffer[!clk]) begin
          $fwrite(f, "Register (5,7) Value: %h\n", PRED5_7_buffer[clk]);
        end
        if (PRED5_8_buffer[clk] != PRED5_8_buffer[!clk]) begin
          $fwrite(f, "Register (5,8) Value: %h\n", PRED5_8_buffer[clk]);
        end
        if (PRED5_9_buffer[clk] != PRED5_9_buffer[!clk]) begin
          $fwrite(f, "Register (5,9) Value: %h\n", PRED5_9_buffer[clk]);
        end
        if (PRED5_10_buffer[clk] != PRED5_10_buffer[!clk]) begin
          $fwrite(f, "Register (5,10) Value: %h\n", PRED5_10_buffer[clk]);
        end
        if (PRED5_11_buffer[clk] != PRED5_11_buffer[!clk]) begin
          $fwrite(f, "Register (5,11) Value: %h\n", PRED5_11_buffer[clk]);
        end
        if (PRED5_12_buffer[clk] != PRED5_12_buffer[!clk]) begin
          $fwrite(f, "Register (5,12) Value: %h\n", PRED5_12_buffer[clk]);
        end
        if (PRED5_13_buffer[clk] != PRED5_13_buffer[!clk]) begin
          $fwrite(f, "Register (5,13) Value: %h\n", PRED5_13_buffer[clk]);
        end
        if (PRED5_14_buffer[clk] != PRED5_14_buffer[!clk]) begin
          $fwrite(f, "Register (5,14) Value: %h\n", PRED5_14_buffer[clk]);
        end
        if (PRED5_15_buffer[clk] != PRED5_15_buffer[!clk]) begin
          $fwrite(f, "Register (5,15) Value: %h\n", PRED5_15_buffer[clk]);
        end
        if (PRED5_16_buffer[clk] != PRED5_16_buffer[!clk]) begin
          $fwrite(f, "Register (5,16) Value: %h\n", PRED5_16_buffer[clk]);
        end
        if (PRED5_17_buffer[clk] != PRED5_17_buffer[!clk]) begin
          $fwrite(f, "Register (5,17) Value: %h\n", PRED5_17_buffer[clk]);
        end
        if (PRED5_18_buffer[clk] != PRED5_18_buffer[!clk]) begin
          $fwrite(f, "Register (5,18) Value: %h\n", PRED5_18_buffer[clk]);
        end
        if (PRED5_19_buffer[clk] != PRED5_19_buffer[!clk]) begin
          $fwrite(f, "Register (5,19) Value: %h\n", PRED5_19_buffer[clk]);
        end
        if (PRED5_20_buffer[clk] != PRED5_20_buffer[!clk]) begin
          $fwrite(f, "Register (5,20) Value: %h\n", PRED5_20_buffer[clk]);
        end
        if (PRED5_21_buffer[clk] != PRED5_21_buffer[!clk]) begin
          $fwrite(f, "Register (5,21) Value: %h\n", PRED5_21_buffer[clk]);
        end
        if (PRED5_22_buffer[clk] != PRED5_22_buffer[!clk]) begin
          $fwrite(f, "Register (5,22) Value: %h\n", PRED5_22_buffer[clk]);
        end
        if (PRED5_23_buffer[clk] != PRED5_23_buffer[!clk]) begin
          $fwrite(f, "Register (5,23) Value: %h\n", PRED5_23_buffer[clk]);
        end
        if (PRED5_24_buffer[clk] != PRED5_24_buffer[!clk]) begin
          $fwrite(f, "Register (5,24) Value: %h\n", PRED5_24_buffer[clk]);
        end
        if (PRED5_25_buffer[clk] != PRED5_25_buffer[!clk]) begin
          $fwrite(f, "Register (5,25) Value: %h\n", PRED5_25_buffer[clk]);
        end
        if (PRED5_26_buffer[clk] != PRED5_26_buffer[!clk]) begin
          $fwrite(f, "Register (5,26) Value: %h\n", PRED5_26_buffer[clk]);
        end
        if (PRED5_27_buffer[clk] != PRED5_27_buffer[!clk]) begin
          $fwrite(f, "Register (5,27) Value: %h\n", PRED5_27_buffer[clk]);
        end
        if (PRED5_28_buffer[clk] != PRED5_28_buffer[!clk]) begin
          $fwrite(f, "Register (5,28) Value: %h\n", PRED5_28_buffer[clk]);
        end
        if (PRED5_29_buffer[clk] != PRED5_29_buffer[!clk]) begin
          $fwrite(f, "Register (5,29) Value: %h\n", PRED5_29_buffer[clk]);
        end
        if (PRED5_30_buffer[clk] != PRED5_30_buffer[!clk]) begin
          $fwrite(f, "Register (5,30) Value: %h\n", PRED5_30_buffer[clk]);
        end
        if (PRED5_31_buffer[clk] != PRED5_31_buffer[!clk]) begin
          $fwrite(f, "Register (5,31) Value: %h\n", PRED5_31_buffer[clk]);
        end
        if (PRED6_0_buffer[clk] != PRED6_0_buffer[!clk]) begin
          $fwrite(f, "Register (6,0) Value: %h\n", PRED6_0_buffer[clk]);
        end
        if (PRED6_1_buffer[clk] != PRED6_1_buffer[!clk]) begin
          $fwrite(f, "Register (6,1) Value: %h\n", PRED6_1_buffer[clk]);
        end
        if (PRED6_2_buffer[clk] != PRED6_2_buffer[!clk]) begin
          $fwrite(f, "Register (6,2) Value: %h\n", PRED6_2_buffer[clk]);
        end
        if (PRED6_3_buffer[clk] != PRED6_3_buffer[!clk]) begin
          $fwrite(f, "Register (6,3) Value: %h\n", PRED6_3_buffer[clk]);
        end
        if (PRED6_4_buffer[clk] != PRED6_4_buffer[!clk]) begin
          $fwrite(f, "Register (6,4) Value: %h\n", PRED6_4_buffer[clk]);
        end
        if (PRED6_5_buffer[clk] != PRED6_5_buffer[!clk]) begin
          $fwrite(f, "Register (6,5) Value: %h\n", PRED6_5_buffer[clk]);
        end
        if (PRED6_6_buffer[clk] != PRED6_6_buffer[!clk]) begin
          $fwrite(f, "Register (6,6) Value: %h\n", PRED6_6_buffer[clk]);
        end
        if (PRED6_7_buffer[clk] != PRED6_7_buffer[!clk]) begin
          $fwrite(f, "Register (6,7) Value: %h\n", PRED6_7_buffer[clk]);
        end
        if (PRED6_8_buffer[clk] != PRED6_8_buffer[!clk]) begin
          $fwrite(f, "Register (6,8) Value: %h\n", PRED6_8_buffer[clk]);
        end
        if (PRED6_9_buffer[clk] != PRED6_9_buffer[!clk]) begin
          $fwrite(f, "Register (6,9) Value: %h\n", PRED6_9_buffer[clk]);
        end
        if (PRED6_10_buffer[clk] != PRED6_10_buffer[!clk]) begin
          $fwrite(f, "Register (6,10) Value: %h\n", PRED6_10_buffer[clk]);
        end
        if (PRED6_11_buffer[clk] != PRED6_11_buffer[!clk]) begin
          $fwrite(f, "Register (6,11) Value: %h\n", PRED6_11_buffer[clk]);
        end
        if (PRED6_12_buffer[clk] != PRED6_12_buffer[!clk]) begin
          $fwrite(f, "Register (6,12) Value: %h\n", PRED6_12_buffer[clk]);
        end
        if (PRED6_13_buffer[clk] != PRED6_13_buffer[!clk]) begin
          $fwrite(f, "Register (6,13) Value: %h\n", PRED6_13_buffer[clk]);
        end
        if (PRED6_14_buffer[clk] != PRED6_14_buffer[!clk]) begin
          $fwrite(f, "Register (6,14) Value: %h\n", PRED6_14_buffer[clk]);
        end
        if (PRED6_15_buffer[clk] != PRED6_15_buffer[!clk]) begin
          $fwrite(f, "Register (6,15) Value: %h\n", PRED6_15_buffer[clk]);
        end
        if (PRED6_16_buffer[clk] != PRED6_16_buffer[!clk]) begin
          $fwrite(f, "Register (6,16) Value: %h\n", PRED6_16_buffer[clk]);
        end
        if (PRED6_17_buffer[clk] != PRED6_17_buffer[!clk]) begin
          $fwrite(f, "Register (6,17) Value: %h\n", PRED6_17_buffer[clk]);
        end
        if (PRED6_18_buffer[clk] != PRED6_18_buffer[!clk]) begin
          $fwrite(f, "Register (6,18) Value: %h\n", PRED6_18_buffer[clk]);
        end
        if (PRED6_19_buffer[clk] != PRED6_19_buffer[!clk]) begin
          $fwrite(f, "Register (6,19) Value: %h\n", PRED6_19_buffer[clk]);
        end
        if (PRED6_20_buffer[clk] != PRED6_20_buffer[!clk]) begin
          $fwrite(f, "Register (6,20) Value: %h\n", PRED6_20_buffer[clk]);
        end
        if (PRED6_21_buffer[clk] != PRED6_21_buffer[!clk]) begin
          $fwrite(f, "Register (6,21) Value: %h\n", PRED6_21_buffer[clk]);
        end
        if (PRED6_22_buffer[clk] != PRED6_22_buffer[!clk]) begin
          $fwrite(f, "Register (6,22) Value: %h\n", PRED6_22_buffer[clk]);
        end
        if (PRED6_23_buffer[clk] != PRED6_23_buffer[!clk]) begin
          $fwrite(f, "Register (6,23) Value: %h\n", PRED6_23_buffer[clk]);
        end
        if (PRED6_24_buffer[clk] != PRED6_24_buffer[!clk]) begin
          $fwrite(f, "Register (6,24) Value: %h\n", PRED6_24_buffer[clk]);
        end
        if (PRED6_25_buffer[clk] != PRED6_25_buffer[!clk]) begin
          $fwrite(f, "Register (6,25) Value: %h\n", PRED6_25_buffer[clk]);
        end
        if (PRED6_26_buffer[clk] != PRED6_26_buffer[!clk]) begin
          $fwrite(f, "Register (6,26) Value: %h\n", PRED6_26_buffer[clk]);
        end
        if (PRED6_27_buffer[clk] != PRED6_27_buffer[!clk]) begin
          $fwrite(f, "Register (6,27) Value: %h\n", PRED6_27_buffer[clk]);
        end
        if (PRED6_28_buffer[clk] != PRED6_28_buffer[!clk]) begin
          $fwrite(f, "Register (6,28) Value: %h\n", PRED6_28_buffer[clk]);
        end
        if (PRED6_29_buffer[clk] != PRED6_29_buffer[!clk]) begin
          $fwrite(f, "Register (6,29) Value: %h\n", PRED6_29_buffer[clk]);
        end
        if (PRED6_30_buffer[clk] != PRED6_30_buffer[!clk]) begin
          $fwrite(f, "Register (6,30) Value: %h\n", PRED6_30_buffer[clk]);
        end
        if (PRED6_31_buffer[clk] != PRED6_31_buffer[!clk]) begin
          $fwrite(f, "Register (6,31) Value: %h\n", PRED6_31_buffer[clk]);
        end
        if (PRED7_0_buffer[clk] != PRED7_0_buffer[!clk]) begin
          $fwrite(f, "Register (7,0) Value: %h\n", PRED7_0_buffer[clk]);
        end
        if (PRED7_1_buffer[clk] != PRED7_1_buffer[!clk]) begin
          $fwrite(f, "Register (7,1) Value: %h\n", PRED7_1_buffer[clk]);
        end
        if (PRED7_2_buffer[clk] != PRED7_2_buffer[!clk]) begin
          $fwrite(f, "Register (7,2) Value: %h\n", PRED7_2_buffer[clk]);
        end
        if (PRED7_3_buffer[clk] != PRED7_3_buffer[!clk]) begin
          $fwrite(f, "Register (7,3) Value: %h\n", PRED7_3_buffer[clk]);
        end
        if (PRED7_4_buffer[clk] != PRED7_4_buffer[!clk]) begin
          $fwrite(f, "Register (7,4) Value: %h\n", PRED7_4_buffer[clk]);
        end
        if (PRED7_5_buffer[clk] != PRED7_5_buffer[!clk]) begin
          $fwrite(f, "Register (7,5) Value: %h\n", PRED7_5_buffer[clk]);
        end
        if (PRED7_6_buffer[clk] != PRED7_6_buffer[!clk]) begin
          $fwrite(f, "Register (7,6) Value: %h\n", PRED7_6_buffer[clk]);
        end
        if (PRED7_7_buffer[clk] != PRED7_7_buffer[!clk]) begin
          $fwrite(f, "Register (7,7) Value: %h\n", PRED7_7_buffer[clk]);
        end
        if (PRED7_8_buffer[clk] != PRED7_8_buffer[!clk]) begin
          $fwrite(f, "Register (7,8) Value: %h\n", PRED7_8_buffer[clk]);
        end
        if (PRED7_9_buffer[clk] != PRED7_9_buffer[!clk]) begin
          $fwrite(f, "Register (7,9) Value: %h\n", PRED7_9_buffer[clk]);
        end
        if (PRED7_10_buffer[clk] != PRED7_10_buffer[!clk]) begin
          $fwrite(f, "Register (7,10) Value: %h\n", PRED7_10_buffer[clk]);
        end
        if (PRED7_11_buffer[clk] != PRED7_11_buffer[!clk]) begin
          $fwrite(f, "Register (7,11) Value: %h\n", PRED7_11_buffer[clk]);
        end
        if (PRED7_12_buffer[clk] != PRED7_12_buffer[!clk]) begin
          $fwrite(f, "Register (7,12) Value: %h\n", PRED7_12_buffer[clk]);
        end
        if (PRED7_13_buffer[clk] != PRED7_13_buffer[!clk]) begin
          $fwrite(f, "Register (7,13) Value: %h\n", PRED7_13_buffer[clk]);
        end
        if (PRED7_14_buffer[clk] != PRED7_14_buffer[!clk]) begin
          $fwrite(f, "Register (7,14) Value: %h\n", PRED7_14_buffer[clk]);
        end
        if (PRED7_15_buffer[clk] != PRED7_15_buffer[!clk]) begin
          $fwrite(f, "Register (7,15) Value: %h\n", PRED7_15_buffer[clk]);
        end
        if (PRED7_16_buffer[clk] != PRED7_16_buffer[!clk]) begin
          $fwrite(f, "Register (7,16) Value: %h\n", PRED7_16_buffer[clk]);
        end
        if (PRED7_17_buffer[clk] != PRED7_17_buffer[!clk]) begin
          $fwrite(f, "Register (7,17) Value: %h\n", PRED7_17_buffer[clk]);
        end
        if (PRED7_18_buffer[clk] != PRED7_18_buffer[!clk]) begin
          $fwrite(f, "Register (7,18) Value: %h\n", PRED7_18_buffer[clk]);
        end
        if (PRED7_19_buffer[clk] != PRED7_19_buffer[!clk]) begin
          $fwrite(f, "Register (7,19) Value: %h\n", PRED7_19_buffer[clk]);
        end
        if (PRED7_20_buffer[clk] != PRED7_20_buffer[!clk]) begin
          $fwrite(f, "Register (7,20) Value: %h\n", PRED7_20_buffer[clk]);
        end
        if (PRED7_21_buffer[clk] != PRED7_21_buffer[!clk]) begin
          $fwrite(f, "Register (7,21) Value: %h\n", PRED7_21_buffer[clk]);
        end
        if (PRED7_22_buffer[clk] != PRED7_22_buffer[!clk]) begin
          $fwrite(f, "Register (7,22) Value: %h\n", PRED7_22_buffer[clk]);
        end
        if (PRED7_23_buffer[clk] != PRED7_23_buffer[!clk]) begin
          $fwrite(f, "Register (7,23) Value: %h\n", PRED7_23_buffer[clk]);
        end
        if (PRED7_24_buffer[clk] != PRED7_24_buffer[!clk]) begin
          $fwrite(f, "Register (7,24) Value: %h\n", PRED7_24_buffer[clk]);
        end
        if (PRED7_25_buffer[clk] != PRED7_25_buffer[!clk]) begin
          $fwrite(f, "Register (7,25) Value: %h\n", PRED7_25_buffer[clk]);
        end
        if (PRED7_26_buffer[clk] != PRED7_26_buffer[!clk]) begin
          $fwrite(f, "Register (7,26) Value: %h\n", PRED7_26_buffer[clk]);
        end
        if (PRED7_27_buffer[clk] != PRED7_27_buffer[!clk]) begin
          $fwrite(f, "Register (7,27) Value: %h\n", PRED7_27_buffer[clk]);
        end
        if (PRED7_28_buffer[clk] != PRED7_28_buffer[!clk]) begin
          $fwrite(f, "Register (7,28) Value: %h\n", PRED7_28_buffer[clk]);
        end
        if (PRED7_29_buffer[clk] != PRED7_29_buffer[!clk]) begin
          $fwrite(f, "Register (7,29) Value: %h\n", PRED7_29_buffer[clk]);
        end
        if (PRED7_30_buffer[clk] != PRED7_30_buffer[!clk]) begin
          $fwrite(f, "Register (7,30) Value: %h\n", PRED7_30_buffer[clk]);
        end
        if (PRED7_31_buffer[clk] != PRED7_31_buffer[!clk]) begin
          $fwrite(f, "Register (7,31) Value: %h\n", PRED7_31_buffer[clk]);
        end
        if (PRED8_0_buffer[clk] != PRED8_0_buffer[!clk]) begin
          $fwrite(f, "Register (8,0) Value: %h\n", PRED8_0_buffer[clk]);
        end
        if (PRED8_1_buffer[clk] != PRED8_1_buffer[!clk]) begin
          $fwrite(f, "Register (8,1) Value: %h\n", PRED8_1_buffer[clk]);
        end
        if (PRED8_2_buffer[clk] != PRED8_2_buffer[!clk]) begin
          $fwrite(f, "Register (8,2) Value: %h\n", PRED8_2_buffer[clk]);
        end
        if (PRED8_3_buffer[clk] != PRED8_3_buffer[!clk]) begin
          $fwrite(f, "Register (8,3) Value: %h\n", PRED8_3_buffer[clk]);
        end
        if (PRED8_4_buffer[clk] != PRED8_4_buffer[!clk]) begin
          $fwrite(f, "Register (8,4) Value: %h\n", PRED8_4_buffer[clk]);
        end
        if (PRED8_5_buffer[clk] != PRED8_5_buffer[!clk]) begin
          $fwrite(f, "Register (8,5) Value: %h\n", PRED8_5_buffer[clk]);
        end
        if (PRED8_6_buffer[clk] != PRED8_6_buffer[!clk]) begin
          $fwrite(f, "Register (8,6) Value: %h\n", PRED8_6_buffer[clk]);
        end
        if (PRED8_7_buffer[clk] != PRED8_7_buffer[!clk]) begin
          $fwrite(f, "Register (8,7) Value: %h\n", PRED8_7_buffer[clk]);
        end
        if (PRED8_8_buffer[clk] != PRED8_8_buffer[!clk]) begin
          $fwrite(f, "Register (8,8) Value: %h\n", PRED8_8_buffer[clk]);
        end
        if (PRED8_9_buffer[clk] != PRED8_9_buffer[!clk]) begin
          $fwrite(f, "Register (8,9) Value: %h\n", PRED8_9_buffer[clk]);
        end
        if (PRED8_10_buffer[clk] != PRED8_10_buffer[!clk]) begin
          $fwrite(f, "Register (8,10) Value: %h\n", PRED8_10_buffer[clk]);
        end
        if (PRED8_11_buffer[clk] != PRED8_11_buffer[!clk]) begin
          $fwrite(f, "Register (8,11) Value: %h\n", PRED8_11_buffer[clk]);
        end
        if (PRED8_12_buffer[clk] != PRED8_12_buffer[!clk]) begin
          $fwrite(f, "Register (8,12) Value: %h\n", PRED8_12_buffer[clk]);
        end
        if (PRED8_13_buffer[clk] != PRED8_13_buffer[!clk]) begin
          $fwrite(f, "Register (8,13) Value: %h\n", PRED8_13_buffer[clk]);
        end
        if (PRED8_14_buffer[clk] != PRED8_14_buffer[!clk]) begin
          $fwrite(f, "Register (8,14) Value: %h\n", PRED8_14_buffer[clk]);
        end
        if (PRED8_15_buffer[clk] != PRED8_15_buffer[!clk]) begin
          $fwrite(f, "Register (8,15) Value: %h\n", PRED8_15_buffer[clk]);
        end
        if (PRED8_16_buffer[clk] != PRED8_16_buffer[!clk]) begin
          $fwrite(f, "Register (8,16) Value: %h\n", PRED8_16_buffer[clk]);
        end
        if (PRED8_17_buffer[clk] != PRED8_17_buffer[!clk]) begin
          $fwrite(f, "Register (8,17) Value: %h\n", PRED8_17_buffer[clk]);
        end
        if (PRED8_18_buffer[clk] != PRED8_18_buffer[!clk]) begin
          $fwrite(f, "Register (8,18) Value: %h\n", PRED8_18_buffer[clk]);
        end
        if (PRED8_19_buffer[clk] != PRED8_19_buffer[!clk]) begin
          $fwrite(f, "Register (8,19) Value: %h\n", PRED8_19_buffer[clk]);
        end
        if (PRED8_20_buffer[clk] != PRED8_20_buffer[!clk]) begin
          $fwrite(f, "Register (8,20) Value: %h\n", PRED8_20_buffer[clk]);
        end
        if (PRED8_21_buffer[clk] != PRED8_21_buffer[!clk]) begin
          $fwrite(f, "Register (8,21) Value: %h\n", PRED8_21_buffer[clk]);
        end
        if (PRED8_22_buffer[clk] != PRED8_22_buffer[!clk]) begin
          $fwrite(f, "Register (8,22) Value: %h\n", PRED8_22_buffer[clk]);
        end
        if (PRED8_23_buffer[clk] != PRED8_23_buffer[!clk]) begin
          $fwrite(f, "Register (8,23) Value: %h\n", PRED8_23_buffer[clk]);
        end
        if (PRED8_24_buffer[clk] != PRED8_24_buffer[!clk]) begin
          $fwrite(f, "Register (8,24) Value: %h\n", PRED8_24_buffer[clk]);
        end
        if (PRED8_25_buffer[clk] != PRED8_25_buffer[!clk]) begin
          $fwrite(f, "Register (8,25) Value: %h\n", PRED8_25_buffer[clk]);
        end
        if (PRED8_26_buffer[clk] != PRED8_26_buffer[!clk]) begin
          $fwrite(f, "Register (8,26) Value: %h\n", PRED8_26_buffer[clk]);
        end
        if (PRED8_27_buffer[clk] != PRED8_27_buffer[!clk]) begin
          $fwrite(f, "Register (8,27) Value: %h\n", PRED8_27_buffer[clk]);
        end
        if (PRED8_28_buffer[clk] != PRED8_28_buffer[!clk]) begin
          $fwrite(f, "Register (8,28) Value: %h\n", PRED8_28_buffer[clk]);
        end
        if (PRED8_29_buffer[clk] != PRED8_29_buffer[!clk]) begin
          $fwrite(f, "Register (8,29) Value: %h\n", PRED8_29_buffer[clk]);
        end
        if (PRED8_30_buffer[clk] != PRED8_30_buffer[!clk]) begin
          $fwrite(f, "Register (8,30) Value: %h\n", PRED8_30_buffer[clk]);
        end
        if (PRED8_31_buffer[clk] != PRED8_31_buffer[!clk]) begin
          $fwrite(f, "Register (8,31) Value: %h\n", PRED8_31_buffer[clk]);
        end
        if (PRED9_0_buffer[clk] != PRED9_0_buffer[!clk]) begin
          $fwrite(f, "Register (9,0) Value: %h\n", PRED9_0_buffer[clk]);
        end
        if (PRED9_1_buffer[clk] != PRED9_1_buffer[!clk]) begin
          $fwrite(f, "Register (9,1) Value: %h\n", PRED9_1_buffer[clk]);
        end
        if (PRED9_2_buffer[clk] != PRED9_2_buffer[!clk]) begin
          $fwrite(f, "Register (9,2) Value: %h\n", PRED9_2_buffer[clk]);
        end
        if (PRED9_3_buffer[clk] != PRED9_3_buffer[!clk]) begin
          $fwrite(f, "Register (9,3) Value: %h\n", PRED9_3_buffer[clk]);
        end
        if (PRED9_4_buffer[clk] != PRED9_4_buffer[!clk]) begin
          $fwrite(f, "Register (9,4) Value: %h\n", PRED9_4_buffer[clk]);
        end
        if (PRED9_5_buffer[clk] != PRED9_5_buffer[!clk]) begin
          $fwrite(f, "Register (9,5) Value: %h\n", PRED9_5_buffer[clk]);
        end
        if (PRED9_6_buffer[clk] != PRED9_6_buffer[!clk]) begin
          $fwrite(f, "Register (9,6) Value: %h\n", PRED9_6_buffer[clk]);
        end
        if (PRED9_7_buffer[clk] != PRED9_7_buffer[!clk]) begin
          $fwrite(f, "Register (9,7) Value: %h\n", PRED9_7_buffer[clk]);
        end
        if (PRED9_8_buffer[clk] != PRED9_8_buffer[!clk]) begin
          $fwrite(f, "Register (9,8) Value: %h\n", PRED9_8_buffer[clk]);
        end
        if (PRED9_9_buffer[clk] != PRED9_9_buffer[!clk]) begin
          $fwrite(f, "Register (9,9) Value: %h\n", PRED9_9_buffer[clk]);
        end
        if (PRED9_10_buffer[clk] != PRED9_10_buffer[!clk]) begin
          $fwrite(f, "Register (9,10) Value: %h\n", PRED9_10_buffer[clk]);
        end
        if (PRED9_11_buffer[clk] != PRED9_11_buffer[!clk]) begin
          $fwrite(f, "Register (9,11) Value: %h\n", PRED9_11_buffer[clk]);
        end
        if (PRED9_12_buffer[clk] != PRED9_12_buffer[!clk]) begin
          $fwrite(f, "Register (9,12) Value: %h\n", PRED9_12_buffer[clk]);
        end
        if (PRED9_13_buffer[clk] != PRED9_13_buffer[!clk]) begin
          $fwrite(f, "Register (9,13) Value: %h\n", PRED9_13_buffer[clk]);
        end
        if (PRED9_14_buffer[clk] != PRED9_14_buffer[!clk]) begin
          $fwrite(f, "Register (9,14) Value: %h\n", PRED9_14_buffer[clk]);
        end
        if (PRED9_15_buffer[clk] != PRED9_15_buffer[!clk]) begin
          $fwrite(f, "Register (9,15) Value: %h\n", PRED9_15_buffer[clk]);
        end
        if (PRED9_16_buffer[clk] != PRED9_16_buffer[!clk]) begin
          $fwrite(f, "Register (9,16) Value: %h\n", PRED9_16_buffer[clk]);
        end
        if (PRED9_17_buffer[clk] != PRED9_17_buffer[!clk]) begin
          $fwrite(f, "Register (9,17) Value: %h\n", PRED9_17_buffer[clk]);
        end
        if (PRED9_18_buffer[clk] != PRED9_18_buffer[!clk]) begin
          $fwrite(f, "Register (9,18) Value: %h\n", PRED9_18_buffer[clk]);
        end
        if (PRED9_19_buffer[clk] != PRED9_19_buffer[!clk]) begin
          $fwrite(f, "Register (9,19) Value: %h\n", PRED9_19_buffer[clk]);
        end
        if (PRED9_20_buffer[clk] != PRED9_20_buffer[!clk]) begin
          $fwrite(f, "Register (9,20) Value: %h\n", PRED9_20_buffer[clk]);
        end
        if (PRED9_21_buffer[clk] != PRED9_21_buffer[!clk]) begin
          $fwrite(f, "Register (9,21) Value: %h\n", PRED9_21_buffer[clk]);
        end
        if (PRED9_22_buffer[clk] != PRED9_22_buffer[!clk]) begin
          $fwrite(f, "Register (9,22) Value: %h\n", PRED9_22_buffer[clk]);
        end
        if (PRED9_23_buffer[clk] != PRED9_23_buffer[!clk]) begin
          $fwrite(f, "Register (9,23) Value: %h\n", PRED9_23_buffer[clk]);
        end
        if (PRED9_24_buffer[clk] != PRED9_24_buffer[!clk]) begin
          $fwrite(f, "Register (9,24) Value: %h\n", PRED9_24_buffer[clk]);
        end
        if (PRED9_25_buffer[clk] != PRED9_25_buffer[!clk]) begin
          $fwrite(f, "Register (9,25) Value: %h\n", PRED9_25_buffer[clk]);
        end
        if (PRED9_26_buffer[clk] != PRED9_26_buffer[!clk]) begin
          $fwrite(f, "Register (9,26) Value: %h\n", PRED9_26_buffer[clk]);
        end
        if (PRED9_27_buffer[clk] != PRED9_27_buffer[!clk]) begin
          $fwrite(f, "Register (9,27) Value: %h\n", PRED9_27_buffer[clk]);
        end
        if (PRED9_28_buffer[clk] != PRED9_28_buffer[!clk]) begin
          $fwrite(f, "Register (9,28) Value: %h\n", PRED9_28_buffer[clk]);
        end
        if (PRED9_29_buffer[clk] != PRED9_29_buffer[!clk]) begin
          $fwrite(f, "Register (9,29) Value: %h\n", PRED9_29_buffer[clk]);
        end
        if (PRED9_30_buffer[clk] != PRED9_30_buffer[!clk]) begin
          $fwrite(f, "Register (9,30) Value: %h\n", PRED9_30_buffer[clk]);
        end
        if (PRED9_31_buffer[clk] != PRED9_31_buffer[!clk]) begin
          $fwrite(f, "Register (9,31) Value: %h\n", PRED9_31_buffer[clk]);
        end
        if (PRED10_0_buffer[clk] != PRED10_0_buffer[!clk]) begin
          $fwrite(f, "Register (10,0) Value: %h\n", PRED10_0_buffer[clk]);
        end
        if (PRED10_1_buffer[clk] != PRED10_1_buffer[!clk]) begin
          $fwrite(f, "Register (10,1) Value: %h\n", PRED10_1_buffer[clk]);
        end
        if (PRED10_2_buffer[clk] != PRED10_2_buffer[!clk]) begin
          $fwrite(f, "Register (10,2) Value: %h\n", PRED10_2_buffer[clk]);
        end
        if (PRED10_3_buffer[clk] != PRED10_3_buffer[!clk]) begin
          $fwrite(f, "Register (10,3) Value: %h\n", PRED10_3_buffer[clk]);
        end
        if (PRED10_4_buffer[clk] != PRED10_4_buffer[!clk]) begin
          $fwrite(f, "Register (10,4) Value: %h\n", PRED10_4_buffer[clk]);
        end
        if (PRED10_5_buffer[clk] != PRED10_5_buffer[!clk]) begin
          $fwrite(f, "Register (10,5) Value: %h\n", PRED10_5_buffer[clk]);
        end
        if (PRED10_6_buffer[clk] != PRED10_6_buffer[!clk]) begin
          $fwrite(f, "Register (10,6) Value: %h\n", PRED10_6_buffer[clk]);
        end
        if (PRED10_7_buffer[clk] != PRED10_7_buffer[!clk]) begin
          $fwrite(f, "Register (10,7) Value: %h\n", PRED10_7_buffer[clk]);
        end
        if (PRED10_8_buffer[clk] != PRED10_8_buffer[!clk]) begin
          $fwrite(f, "Register (10,8) Value: %h\n", PRED10_8_buffer[clk]);
        end
        if (PRED10_9_buffer[clk] != PRED10_9_buffer[!clk]) begin
          $fwrite(f, "Register (10,9) Value: %h\n", PRED10_9_buffer[clk]);
        end
        if (PRED10_10_buffer[clk] != PRED10_10_buffer[!clk]) begin
          $fwrite(f, "Register (10,10) Value: %h\n", PRED10_10_buffer[clk]);
        end
        if (PRED10_11_buffer[clk] != PRED10_11_buffer[!clk]) begin
          $fwrite(f, "Register (10,11) Value: %h\n", PRED10_11_buffer[clk]);
        end
        if (PRED10_12_buffer[clk] != PRED10_12_buffer[!clk]) begin
          $fwrite(f, "Register (10,12) Value: %h\n", PRED10_12_buffer[clk]);
        end
        if (PRED10_13_buffer[clk] != PRED10_13_buffer[!clk]) begin
          $fwrite(f, "Register (10,13) Value: %h\n", PRED10_13_buffer[clk]);
        end
        if (PRED10_14_buffer[clk] != PRED10_14_buffer[!clk]) begin
          $fwrite(f, "Register (10,14) Value: %h\n", PRED10_14_buffer[clk]);
        end
        if (PRED10_15_buffer[clk] != PRED10_15_buffer[!clk]) begin
          $fwrite(f, "Register (10,15) Value: %h\n", PRED10_15_buffer[clk]);
        end
        if (PRED10_16_buffer[clk] != PRED10_16_buffer[!clk]) begin
          $fwrite(f, "Register (10,16) Value: %h\n", PRED10_16_buffer[clk]);
        end
        if (PRED10_17_buffer[clk] != PRED10_17_buffer[!clk]) begin
          $fwrite(f, "Register (10,17) Value: %h\n", PRED10_17_buffer[clk]);
        end
        if (PRED10_18_buffer[clk] != PRED10_18_buffer[!clk]) begin
          $fwrite(f, "Register (10,18) Value: %h\n", PRED10_18_buffer[clk]);
        end
        if (PRED10_19_buffer[clk] != PRED10_19_buffer[!clk]) begin
          $fwrite(f, "Register (10,19) Value: %h\n", PRED10_19_buffer[clk]);
        end
        if (PRED10_20_buffer[clk] != PRED10_20_buffer[!clk]) begin
          $fwrite(f, "Register (10,20) Value: %h\n", PRED10_20_buffer[clk]);
        end
        if (PRED10_21_buffer[clk] != PRED10_21_buffer[!clk]) begin
          $fwrite(f, "Register (10,21) Value: %h\n", PRED10_21_buffer[clk]);
        end
        if (PRED10_22_buffer[clk] != PRED10_22_buffer[!clk]) begin
          $fwrite(f, "Register (10,22) Value: %h\n", PRED10_22_buffer[clk]);
        end
        if (PRED10_23_buffer[clk] != PRED10_23_buffer[!clk]) begin
          $fwrite(f, "Register (10,23) Value: %h\n", PRED10_23_buffer[clk]);
        end
        if (PRED10_24_buffer[clk] != PRED10_24_buffer[!clk]) begin
          $fwrite(f, "Register (10,24) Value: %h\n", PRED10_24_buffer[clk]);
        end
        if (PRED10_25_buffer[clk] != PRED10_25_buffer[!clk]) begin
          $fwrite(f, "Register (10,25) Value: %h\n", PRED10_25_buffer[clk]);
        end
        if (PRED10_26_buffer[clk] != PRED10_26_buffer[!clk]) begin
          $fwrite(f, "Register (10,26) Value: %h\n", PRED10_26_buffer[clk]);
        end
        if (PRED10_27_buffer[clk] != PRED10_27_buffer[!clk]) begin
          $fwrite(f, "Register (10,27) Value: %h\n", PRED10_27_buffer[clk]);
        end
        if (PRED10_28_buffer[clk] != PRED10_28_buffer[!clk]) begin
          $fwrite(f, "Register (10,28) Value: %h\n", PRED10_28_buffer[clk]);
        end
        if (PRED10_29_buffer[clk] != PRED10_29_buffer[!clk]) begin
          $fwrite(f, "Register (10,29) Value: %h\n", PRED10_29_buffer[clk]);
        end
        if (PRED10_30_buffer[clk] != PRED10_30_buffer[!clk]) begin
          $fwrite(f, "Register (10,30) Value: %h\n", PRED10_30_buffer[clk]);
        end
        if (PRED10_31_buffer[clk] != PRED10_31_buffer[!clk]) begin
          $fwrite(f, "Register (10,31) Value: %h\n", PRED10_31_buffer[clk]);
        end
        if (PRED11_0_buffer[clk] != PRED11_0_buffer[!clk]) begin
          $fwrite(f, "Register (11,0) Value: %h\n", PRED11_0_buffer[clk]);
        end
        if (PRED11_1_buffer[clk] != PRED11_1_buffer[!clk]) begin
          $fwrite(f, "Register (11,1) Value: %h\n", PRED11_1_buffer[clk]);
        end
        if (PRED11_2_buffer[clk] != PRED11_2_buffer[!clk]) begin
          $fwrite(f, "Register (11,2) Value: %h\n", PRED11_2_buffer[clk]);
        end
        if (PRED11_3_buffer[clk] != PRED11_3_buffer[!clk]) begin
          $fwrite(f, "Register (11,3) Value: %h\n", PRED11_3_buffer[clk]);
        end
        if (PRED11_4_buffer[clk] != PRED11_4_buffer[!clk]) begin
          $fwrite(f, "Register (11,4) Value: %h\n", PRED11_4_buffer[clk]);
        end
        if (PRED11_5_buffer[clk] != PRED11_5_buffer[!clk]) begin
          $fwrite(f, "Register (11,5) Value: %h\n", PRED11_5_buffer[clk]);
        end
        if (PRED11_6_buffer[clk] != PRED11_6_buffer[!clk]) begin
          $fwrite(f, "Register (11,6) Value: %h\n", PRED11_6_buffer[clk]);
        end
        if (PRED11_7_buffer[clk] != PRED11_7_buffer[!clk]) begin
          $fwrite(f, "Register (11,7) Value: %h\n", PRED11_7_buffer[clk]);
        end
        if (PRED11_8_buffer[clk] != PRED11_8_buffer[!clk]) begin
          $fwrite(f, "Register (11,8) Value: %h\n", PRED11_8_buffer[clk]);
        end
        if (PRED11_9_buffer[clk] != PRED11_9_buffer[!clk]) begin
          $fwrite(f, "Register (11,9) Value: %h\n", PRED11_9_buffer[clk]);
        end
        if (PRED11_10_buffer[clk] != PRED11_10_buffer[!clk]) begin
          $fwrite(f, "Register (11,10) Value: %h\n", PRED11_10_buffer[clk]);
        end
        if (PRED11_11_buffer[clk] != PRED11_11_buffer[!clk]) begin
          $fwrite(f, "Register (11,11) Value: %h\n", PRED11_11_buffer[clk]);
        end
        if (PRED11_12_buffer[clk] != PRED11_12_buffer[!clk]) begin
          $fwrite(f, "Register (11,12) Value: %h\n", PRED11_12_buffer[clk]);
        end
        if (PRED11_13_buffer[clk] != PRED11_13_buffer[!clk]) begin
          $fwrite(f, "Register (11,13) Value: %h\n", PRED11_13_buffer[clk]);
        end
        if (PRED11_14_buffer[clk] != PRED11_14_buffer[!clk]) begin
          $fwrite(f, "Register (11,14) Value: %h\n", PRED11_14_buffer[clk]);
        end
        if (PRED11_15_buffer[clk] != PRED11_15_buffer[!clk]) begin
          $fwrite(f, "Register (11,15) Value: %h\n", PRED11_15_buffer[clk]);
        end
        if (PRED11_16_buffer[clk] != PRED11_16_buffer[!clk]) begin
          $fwrite(f, "Register (11,16) Value: %h\n", PRED11_16_buffer[clk]);
        end
        if (PRED11_17_buffer[clk] != PRED11_17_buffer[!clk]) begin
          $fwrite(f, "Register (11,17) Value: %h\n", PRED11_17_buffer[clk]);
        end
        if (PRED11_18_buffer[clk] != PRED11_18_buffer[!clk]) begin
          $fwrite(f, "Register (11,18) Value: %h\n", PRED11_18_buffer[clk]);
        end
        if (PRED11_19_buffer[clk] != PRED11_19_buffer[!clk]) begin
          $fwrite(f, "Register (11,19) Value: %h\n", PRED11_19_buffer[clk]);
        end
        if (PRED11_20_buffer[clk] != PRED11_20_buffer[!clk]) begin
          $fwrite(f, "Register (11,20) Value: %h\n", PRED11_20_buffer[clk]);
        end
        if (PRED11_21_buffer[clk] != PRED11_21_buffer[!clk]) begin
          $fwrite(f, "Register (11,21) Value: %h\n", PRED11_21_buffer[clk]);
        end
        if (PRED11_22_buffer[clk] != PRED11_22_buffer[!clk]) begin
          $fwrite(f, "Register (11,22) Value: %h\n", PRED11_22_buffer[clk]);
        end
        if (PRED11_23_buffer[clk] != PRED11_23_buffer[!clk]) begin
          $fwrite(f, "Register (11,23) Value: %h\n", PRED11_23_buffer[clk]);
        end
        if (PRED11_24_buffer[clk] != PRED11_24_buffer[!clk]) begin
          $fwrite(f, "Register (11,24) Value: %h\n", PRED11_24_buffer[clk]);
        end
        if (PRED11_25_buffer[clk] != PRED11_25_buffer[!clk]) begin
          $fwrite(f, "Register (11,25) Value: %h\n", PRED11_25_buffer[clk]);
        end
        if (PRED11_26_buffer[clk] != PRED11_26_buffer[!clk]) begin
          $fwrite(f, "Register (11,26) Value: %h\n", PRED11_26_buffer[clk]);
        end
        if (PRED11_27_buffer[clk] != PRED11_27_buffer[!clk]) begin
          $fwrite(f, "Register (11,27) Value: %h\n", PRED11_27_buffer[clk]);
        end
        if (PRED11_28_buffer[clk] != PRED11_28_buffer[!clk]) begin
          $fwrite(f, "Register (11,28) Value: %h\n", PRED11_28_buffer[clk]);
        end
        if (PRED11_29_buffer[clk] != PRED11_29_buffer[!clk]) begin
          $fwrite(f, "Register (11,29) Value: %h\n", PRED11_29_buffer[clk]);
        end
        if (PRED11_30_buffer[clk] != PRED11_30_buffer[!clk]) begin
          $fwrite(f, "Register (11,30) Value: %h\n", PRED11_30_buffer[clk]);
        end
        if (PRED11_31_buffer[clk] != PRED11_31_buffer[!clk]) begin
          $fwrite(f, "Register (11,31) Value: %h\n", PRED11_31_buffer[clk]);
        end
        if (PRED12_0_buffer[clk] != PRED12_0_buffer[!clk]) begin
          $fwrite(f, "Register (12,0) Value: %h\n", PRED12_0_buffer[clk]);
        end
        if (PRED12_1_buffer[clk] != PRED12_1_buffer[!clk]) begin
          $fwrite(f, "Register (12,1) Value: %h\n", PRED12_1_buffer[clk]);
        end
        if (PRED12_2_buffer[clk] != PRED12_2_buffer[!clk]) begin
          $fwrite(f, "Register (12,2) Value: %h\n", PRED12_2_buffer[clk]);
        end
        if (PRED12_3_buffer[clk] != PRED12_3_buffer[!clk]) begin
          $fwrite(f, "Register (12,3) Value: %h\n", PRED12_3_buffer[clk]);
        end
        if (PRED12_4_buffer[clk] != PRED12_4_buffer[!clk]) begin
          $fwrite(f, "Register (12,4) Value: %h\n", PRED12_4_buffer[clk]);
        end
        if (PRED12_5_buffer[clk] != PRED12_5_buffer[!clk]) begin
          $fwrite(f, "Register (12,5) Value: %h\n", PRED12_5_buffer[clk]);
        end
        if (PRED12_6_buffer[clk] != PRED12_6_buffer[!clk]) begin
          $fwrite(f, "Register (12,6) Value: %h\n", PRED12_6_buffer[clk]);
        end
        if (PRED12_7_buffer[clk] != PRED12_7_buffer[!clk]) begin
          $fwrite(f, "Register (12,7) Value: %h\n", PRED12_7_buffer[clk]);
        end
        if (PRED12_8_buffer[clk] != PRED12_8_buffer[!clk]) begin
          $fwrite(f, "Register (12,8) Value: %h\n", PRED12_8_buffer[clk]);
        end
        if (PRED12_9_buffer[clk] != PRED12_9_buffer[!clk]) begin
          $fwrite(f, "Register (12,9) Value: %h\n", PRED12_9_buffer[clk]);
        end
        if (PRED12_10_buffer[clk] != PRED12_10_buffer[!clk]) begin
          $fwrite(f, "Register (12,10) Value: %h\n", PRED12_10_buffer[clk]);
        end
        if (PRED12_11_buffer[clk] != PRED12_11_buffer[!clk]) begin
          $fwrite(f, "Register (12,11) Value: %h\n", PRED12_11_buffer[clk]);
        end
        if (PRED12_12_buffer[clk] != PRED12_12_buffer[!clk]) begin
          $fwrite(f, "Register (12,12) Value: %h\n", PRED12_12_buffer[clk]);
        end
        if (PRED12_13_buffer[clk] != PRED12_13_buffer[!clk]) begin
          $fwrite(f, "Register (12,13) Value: %h\n", PRED12_13_buffer[clk]);
        end
        if (PRED12_14_buffer[clk] != PRED12_14_buffer[!clk]) begin
          $fwrite(f, "Register (12,14) Value: %h\n", PRED12_14_buffer[clk]);
        end
        if (PRED12_15_buffer[clk] != PRED12_15_buffer[!clk]) begin
          $fwrite(f, "Register (12,15) Value: %h\n", PRED12_15_buffer[clk]);
        end
        if (PRED12_16_buffer[clk] != PRED12_16_buffer[!clk]) begin
          $fwrite(f, "Register (12,16) Value: %h\n", PRED12_16_buffer[clk]);
        end
        if (PRED12_17_buffer[clk] != PRED12_17_buffer[!clk]) begin
          $fwrite(f, "Register (12,17) Value: %h\n", PRED12_17_buffer[clk]);
        end
        if (PRED12_18_buffer[clk] != PRED12_18_buffer[!clk]) begin
          $fwrite(f, "Register (12,18) Value: %h\n", PRED12_18_buffer[clk]);
        end
        if (PRED12_19_buffer[clk] != PRED12_19_buffer[!clk]) begin
          $fwrite(f, "Register (12,19) Value: %h\n", PRED12_19_buffer[clk]);
        end
        if (PRED12_20_buffer[clk] != PRED12_20_buffer[!clk]) begin
          $fwrite(f, "Register (12,20) Value: %h\n", PRED12_20_buffer[clk]);
        end
        if (PRED12_21_buffer[clk] != PRED12_21_buffer[!clk]) begin
          $fwrite(f, "Register (12,21) Value: %h\n", PRED12_21_buffer[clk]);
        end
        if (PRED12_22_buffer[clk] != PRED12_22_buffer[!clk]) begin
          $fwrite(f, "Register (12,22) Value: %h\n", PRED12_22_buffer[clk]);
        end
        if (PRED12_23_buffer[clk] != PRED12_23_buffer[!clk]) begin
          $fwrite(f, "Register (12,23) Value: %h\n", PRED12_23_buffer[clk]);
        end
        if (PRED12_24_buffer[clk] != PRED12_24_buffer[!clk]) begin
          $fwrite(f, "Register (12,24) Value: %h\n", PRED12_24_buffer[clk]);
        end
        if (PRED12_25_buffer[clk] != PRED12_25_buffer[!clk]) begin
          $fwrite(f, "Register (12,25) Value: %h\n", PRED12_25_buffer[clk]);
        end
        if (PRED12_26_buffer[clk] != PRED12_26_buffer[!clk]) begin
          $fwrite(f, "Register (12,26) Value: %h\n", PRED12_26_buffer[clk]);
        end
        if (PRED12_27_buffer[clk] != PRED12_27_buffer[!clk]) begin
          $fwrite(f, "Register (12,27) Value: %h\n", PRED12_27_buffer[clk]);
        end
        if (PRED12_28_buffer[clk] != PRED12_28_buffer[!clk]) begin
          $fwrite(f, "Register (12,28) Value: %h\n", PRED12_28_buffer[clk]);
        end
        if (PRED12_29_buffer[clk] != PRED12_29_buffer[!clk]) begin
          $fwrite(f, "Register (12,29) Value: %h\n", PRED12_29_buffer[clk]);
        end
        if (PRED12_30_buffer[clk] != PRED12_30_buffer[!clk]) begin
          $fwrite(f, "Register (12,30) Value: %h\n", PRED12_30_buffer[clk]);
        end
        if (PRED12_31_buffer[clk] != PRED12_31_buffer[!clk]) begin
          $fwrite(f, "Register (12,31) Value: %h\n", PRED12_31_buffer[clk]);
        end
        if (PRED13_0_buffer[clk] != PRED13_0_buffer[!clk]) begin
          $fwrite(f, "Register (13,0) Value: %h\n", PRED13_0_buffer[clk]);
        end
        if (PRED13_1_buffer[clk] != PRED13_1_buffer[!clk]) begin
          $fwrite(f, "Register (13,1) Value: %h\n", PRED13_1_buffer[clk]);
        end
        if (PRED13_2_buffer[clk] != PRED13_2_buffer[!clk]) begin
          $fwrite(f, "Register (13,2) Value: %h\n", PRED13_2_buffer[clk]);
        end
        if (PRED13_3_buffer[clk] != PRED13_3_buffer[!clk]) begin
          $fwrite(f, "Register (13,3) Value: %h\n", PRED13_3_buffer[clk]);
        end
        if (PRED13_4_buffer[clk] != PRED13_4_buffer[!clk]) begin
          $fwrite(f, "Register (13,4) Value: %h\n", PRED13_4_buffer[clk]);
        end
        if (PRED13_5_buffer[clk] != PRED13_5_buffer[!clk]) begin
          $fwrite(f, "Register (13,5) Value: %h\n", PRED13_5_buffer[clk]);
        end
        if (PRED13_6_buffer[clk] != PRED13_6_buffer[!clk]) begin
          $fwrite(f, "Register (13,6) Value: %h\n", PRED13_6_buffer[clk]);
        end
        if (PRED13_7_buffer[clk] != PRED13_7_buffer[!clk]) begin
          $fwrite(f, "Register (13,7) Value: %h\n", PRED13_7_buffer[clk]);
        end
        if (PRED13_8_buffer[clk] != PRED13_8_buffer[!clk]) begin
          $fwrite(f, "Register (13,8) Value: %h\n", PRED13_8_buffer[clk]);
        end
        if (PRED13_9_buffer[clk] != PRED13_9_buffer[!clk]) begin
          $fwrite(f, "Register (13,9) Value: %h\n", PRED13_9_buffer[clk]);
        end
        if (PRED13_10_buffer[clk] != PRED13_10_buffer[!clk]) begin
          $fwrite(f, "Register (13,10) Value: %h\n", PRED13_10_buffer[clk]);
        end
        if (PRED13_11_buffer[clk] != PRED13_11_buffer[!clk]) begin
          $fwrite(f, "Register (13,11) Value: %h\n", PRED13_11_buffer[clk]);
        end
        if (PRED13_12_buffer[clk] != PRED13_12_buffer[!clk]) begin
          $fwrite(f, "Register (13,12) Value: %h\n", PRED13_12_buffer[clk]);
        end
        if (PRED13_13_buffer[clk] != PRED13_13_buffer[!clk]) begin
          $fwrite(f, "Register (13,13) Value: %h\n", PRED13_13_buffer[clk]);
        end
        if (PRED13_14_buffer[clk] != PRED13_14_buffer[!clk]) begin
          $fwrite(f, "Register (13,14) Value: %h\n", PRED13_14_buffer[clk]);
        end
        if (PRED13_15_buffer[clk] != PRED13_15_buffer[!clk]) begin
          $fwrite(f, "Register (13,15) Value: %h\n", PRED13_15_buffer[clk]);
        end
        if (PRED13_16_buffer[clk] != PRED13_16_buffer[!clk]) begin
          $fwrite(f, "Register (13,16) Value: %h\n", PRED13_16_buffer[clk]);
        end
        if (PRED13_17_buffer[clk] != PRED13_17_buffer[!clk]) begin
          $fwrite(f, "Register (13,17) Value: %h\n", PRED13_17_buffer[clk]);
        end
        if (PRED13_18_buffer[clk] != PRED13_18_buffer[!clk]) begin
          $fwrite(f, "Register (13,18) Value: %h\n", PRED13_18_buffer[clk]);
        end
        if (PRED13_19_buffer[clk] != PRED13_19_buffer[!clk]) begin
          $fwrite(f, "Register (13,19) Value: %h\n", PRED13_19_buffer[clk]);
        end
        if (PRED13_20_buffer[clk] != PRED13_20_buffer[!clk]) begin
          $fwrite(f, "Register (13,20) Value: %h\n", PRED13_20_buffer[clk]);
        end
        if (PRED13_21_buffer[clk] != PRED13_21_buffer[!clk]) begin
          $fwrite(f, "Register (13,21) Value: %h\n", PRED13_21_buffer[clk]);
        end
        if (PRED13_22_buffer[clk] != PRED13_22_buffer[!clk]) begin
          $fwrite(f, "Register (13,22) Value: %h\n", PRED13_22_buffer[clk]);
        end
        if (PRED13_23_buffer[clk] != PRED13_23_buffer[!clk]) begin
          $fwrite(f, "Register (13,23) Value: %h\n", PRED13_23_buffer[clk]);
        end
        if (PRED13_24_buffer[clk] != PRED13_24_buffer[!clk]) begin
          $fwrite(f, "Register (13,24) Value: %h\n", PRED13_24_buffer[clk]);
        end
        if (PRED13_25_buffer[clk] != PRED13_25_buffer[!clk]) begin
          $fwrite(f, "Register (13,25) Value: %h\n", PRED13_25_buffer[clk]);
        end
        if (PRED13_26_buffer[clk] != PRED13_26_buffer[!clk]) begin
          $fwrite(f, "Register (13,26) Value: %h\n", PRED13_26_buffer[clk]);
        end
        if (PRED13_27_buffer[clk] != PRED13_27_buffer[!clk]) begin
          $fwrite(f, "Register (13,27) Value: %h\n", PRED13_27_buffer[clk]);
        end
        if (PRED13_28_buffer[clk] != PRED13_28_buffer[!clk]) begin
          $fwrite(f, "Register (13,28) Value: %h\n", PRED13_28_buffer[clk]);
        end
        if (PRED13_29_buffer[clk] != PRED13_29_buffer[!clk]) begin
          $fwrite(f, "Register (13,29) Value: %h\n", PRED13_29_buffer[clk]);
        end
        if (PRED13_30_buffer[clk] != PRED13_30_buffer[!clk]) begin
          $fwrite(f, "Register (13,30) Value: %h\n", PRED13_30_buffer[clk]);
        end
        if (PRED13_31_buffer[clk] != PRED13_31_buffer[!clk]) begin
          $fwrite(f, "Register (13,31) Value: %h\n", PRED13_31_buffer[clk]);
        end
        if (PRED14_0_buffer[clk] != PRED14_0_buffer[!clk]) begin
          $fwrite(f, "Register (14,0) Value: %h\n", PRED14_0_buffer[clk]);
        end
        if (PRED14_1_buffer[clk] != PRED14_1_buffer[!clk]) begin
          $fwrite(f, "Register (14,1) Value: %h\n", PRED14_1_buffer[clk]);
        end
        if (PRED14_2_buffer[clk] != PRED14_2_buffer[!clk]) begin
          $fwrite(f, "Register (14,2) Value: %h\n", PRED14_2_buffer[clk]);
        end
        if (PRED14_3_buffer[clk] != PRED14_3_buffer[!clk]) begin
          $fwrite(f, "Register (14,3) Value: %h\n", PRED14_3_buffer[clk]);
        end
        if (PRED14_4_buffer[clk] != PRED14_4_buffer[!clk]) begin
          $fwrite(f, "Register (14,4) Value: %h\n", PRED14_4_buffer[clk]);
        end
        if (PRED14_5_buffer[clk] != PRED14_5_buffer[!clk]) begin
          $fwrite(f, "Register (14,5) Value: %h\n", PRED14_5_buffer[clk]);
        end
        if (PRED14_6_buffer[clk] != PRED14_6_buffer[!clk]) begin
          $fwrite(f, "Register (14,6) Value: %h\n", PRED14_6_buffer[clk]);
        end
        if (PRED14_7_buffer[clk] != PRED14_7_buffer[!clk]) begin
          $fwrite(f, "Register (14,7) Value: %h\n", PRED14_7_buffer[clk]);
        end
        if (PRED14_8_buffer[clk] != PRED14_8_buffer[!clk]) begin
          $fwrite(f, "Register (14,8) Value: %h\n", PRED14_8_buffer[clk]);
        end
        if (PRED14_9_buffer[clk] != PRED14_9_buffer[!clk]) begin
          $fwrite(f, "Register (14,9) Value: %h\n", PRED14_9_buffer[clk]);
        end
        if (PRED14_10_buffer[clk] != PRED14_10_buffer[!clk]) begin
          $fwrite(f, "Register (14,10) Value: %h\n", PRED14_10_buffer[clk]);
        end
        if (PRED14_11_buffer[clk] != PRED14_11_buffer[!clk]) begin
          $fwrite(f, "Register (14,11) Value: %h\n", PRED14_11_buffer[clk]);
        end
        if (PRED14_12_buffer[clk] != PRED14_12_buffer[!clk]) begin
          $fwrite(f, "Register (14,12) Value: %h\n", PRED14_12_buffer[clk]);
        end
        if (PRED14_13_buffer[clk] != PRED14_13_buffer[!clk]) begin
          $fwrite(f, "Register (14,13) Value: %h\n", PRED14_13_buffer[clk]);
        end
        if (PRED14_14_buffer[clk] != PRED14_14_buffer[!clk]) begin
          $fwrite(f, "Register (14,14) Value: %h\n", PRED14_14_buffer[clk]);
        end
        if (PRED14_15_buffer[clk] != PRED14_15_buffer[!clk]) begin
          $fwrite(f, "Register (14,15) Value: %h\n", PRED14_15_buffer[clk]);
        end
        if (PRED14_16_buffer[clk] != PRED14_16_buffer[!clk]) begin
          $fwrite(f, "Register (14,16) Value: %h\n", PRED14_16_buffer[clk]);
        end
        if (PRED14_17_buffer[clk] != PRED14_17_buffer[!clk]) begin
          $fwrite(f, "Register (14,17) Value: %h\n", PRED14_17_buffer[clk]);
        end
        if (PRED14_18_buffer[clk] != PRED14_18_buffer[!clk]) begin
          $fwrite(f, "Register (14,18) Value: %h\n", PRED14_18_buffer[clk]);
        end
        if (PRED14_19_buffer[clk] != PRED14_19_buffer[!clk]) begin
          $fwrite(f, "Register (14,19) Value: %h\n", PRED14_19_buffer[clk]);
        end
        if (PRED14_20_buffer[clk] != PRED14_20_buffer[!clk]) begin
          $fwrite(f, "Register (14,20) Value: %h\n", PRED14_20_buffer[clk]);
        end
        if (PRED14_21_buffer[clk] != PRED14_21_buffer[!clk]) begin
          $fwrite(f, "Register (14,21) Value: %h\n", PRED14_21_buffer[clk]);
        end
        if (PRED14_22_buffer[clk] != PRED14_22_buffer[!clk]) begin
          $fwrite(f, "Register (14,22) Value: %h\n", PRED14_22_buffer[clk]);
        end
        if (PRED14_23_buffer[clk] != PRED14_23_buffer[!clk]) begin
          $fwrite(f, "Register (14,23) Value: %h\n", PRED14_23_buffer[clk]);
        end
        if (PRED14_24_buffer[clk] != PRED14_24_buffer[!clk]) begin
          $fwrite(f, "Register (14,24) Value: %h\n", PRED14_24_buffer[clk]);
        end
        if (PRED14_25_buffer[clk] != PRED14_25_buffer[!clk]) begin
          $fwrite(f, "Register (14,25) Value: %h\n", PRED14_25_buffer[clk]);
        end
        if (PRED14_26_buffer[clk] != PRED14_26_buffer[!clk]) begin
          $fwrite(f, "Register (14,26) Value: %h\n", PRED14_26_buffer[clk]);
        end
        if (PRED14_27_buffer[clk] != PRED14_27_buffer[!clk]) begin
          $fwrite(f, "Register (14,27) Value: %h\n", PRED14_27_buffer[clk]);
        end
        if (PRED14_28_buffer[clk] != PRED14_28_buffer[!clk]) begin
          $fwrite(f, "Register (14,28) Value: %h\n", PRED14_28_buffer[clk]);
        end
        if (PRED14_29_buffer[clk] != PRED14_29_buffer[!clk]) begin
          $fwrite(f, "Register (14,29) Value: %h\n", PRED14_29_buffer[clk]);
        end
        if (PRED14_30_buffer[clk] != PRED14_30_buffer[!clk]) begin
          $fwrite(f, "Register (14,30) Value: %h\n", PRED14_30_buffer[clk]);
        end
        if (PRED14_31_buffer[clk] != PRED14_31_buffer[!clk]) begin
          $fwrite(f, "Register (14,31) Value: %h\n", PRED14_31_buffer[clk]);
        end
        if (PRED15_0_buffer[clk] != PRED15_0_buffer[!clk]) begin
          $fwrite(f, "Register (15,0) Value: %h\n", PRED15_0_buffer[clk]);
        end
        if (PRED15_1_buffer[clk] != PRED15_1_buffer[!clk]) begin
          $fwrite(f, "Register (15,1) Value: %h\n", PRED15_1_buffer[clk]);
        end
        if (PRED15_2_buffer[clk] != PRED15_2_buffer[!clk]) begin
          $fwrite(f, "Register (15,2) Value: %h\n", PRED15_2_buffer[clk]);
        end
        if (PRED15_3_buffer[clk] != PRED15_3_buffer[!clk]) begin
          $fwrite(f, "Register (15,3) Value: %h\n", PRED15_3_buffer[clk]);
        end
        if (PRED15_4_buffer[clk] != PRED15_4_buffer[!clk]) begin
          $fwrite(f, "Register (15,4) Value: %h\n", PRED15_4_buffer[clk]);
        end
        if (PRED15_5_buffer[clk] != PRED15_5_buffer[!clk]) begin
          $fwrite(f, "Register (15,5) Value: %h\n", PRED15_5_buffer[clk]);
        end
        if (PRED15_6_buffer[clk] != PRED15_6_buffer[!clk]) begin
          $fwrite(f, "Register (15,6) Value: %h\n", PRED15_6_buffer[clk]);
        end
        if (PRED15_7_buffer[clk] != PRED15_7_buffer[!clk]) begin
          $fwrite(f, "Register (15,7) Value: %h\n", PRED15_7_buffer[clk]);
        end
        if (PRED15_8_buffer[clk] != PRED15_8_buffer[!clk]) begin
          $fwrite(f, "Register (15,8) Value: %h\n", PRED15_8_buffer[clk]);
        end
        if (PRED15_9_buffer[clk] != PRED15_9_buffer[!clk]) begin
          $fwrite(f, "Register (15,9) Value: %h\n", PRED15_9_buffer[clk]);
        end
        if (PRED15_10_buffer[clk] != PRED15_10_buffer[!clk]) begin
          $fwrite(f, "Register (15,10) Value: %h\n", PRED15_10_buffer[clk]);
        end
        if (PRED15_11_buffer[clk] != PRED15_11_buffer[!clk]) begin
          $fwrite(f, "Register (15,11) Value: %h\n", PRED15_11_buffer[clk]);
        end
        if (PRED15_12_buffer[clk] != PRED15_12_buffer[!clk]) begin
          $fwrite(f, "Register (15,12) Value: %h\n", PRED15_12_buffer[clk]);
        end
        if (PRED15_13_buffer[clk] != PRED15_13_buffer[!clk]) begin
          $fwrite(f, "Register (15,13) Value: %h\n", PRED15_13_buffer[clk]);
        end
        if (PRED15_14_buffer[clk] != PRED15_14_buffer[!clk]) begin
          $fwrite(f, "Register (15,14) Value: %h\n", PRED15_14_buffer[clk]);
        end
        if (PRED15_15_buffer[clk] != PRED15_15_buffer[!clk]) begin
          $fwrite(f, "Register (15,15) Value: %h\n", PRED15_15_buffer[clk]);
        end
        if (PRED15_16_buffer[clk] != PRED15_16_buffer[!clk]) begin
          $fwrite(f, "Register (15,16) Value: %h\n", PRED15_16_buffer[clk]);
        end
        if (PRED15_17_buffer[clk] != PRED15_17_buffer[!clk]) begin
          $fwrite(f, "Register (15,17) Value: %h\n", PRED15_17_buffer[clk]);
        end
        if (PRED15_18_buffer[clk] != PRED15_18_buffer[!clk]) begin
          $fwrite(f, "Register (15,18) Value: %h\n", PRED15_18_buffer[clk]);
        end
        if (PRED15_19_buffer[clk] != PRED15_19_buffer[!clk]) begin
          $fwrite(f, "Register (15,19) Value: %h\n", PRED15_19_buffer[clk]);
        end
        if (PRED15_20_buffer[clk] != PRED15_20_buffer[!clk]) begin
          $fwrite(f, "Register (15,20) Value: %h\n", PRED15_20_buffer[clk]);
        end
        if (PRED15_21_buffer[clk] != PRED15_21_buffer[!clk]) begin
          $fwrite(f, "Register (15,21) Value: %h\n", PRED15_21_buffer[clk]);
        end
        if (PRED15_22_buffer[clk] != PRED15_22_buffer[!clk]) begin
          $fwrite(f, "Register (15,22) Value: %h\n", PRED15_22_buffer[clk]);
        end
        if (PRED15_23_buffer[clk] != PRED15_23_buffer[!clk]) begin
          $fwrite(f, "Register (15,23) Value: %h\n", PRED15_23_buffer[clk]);
        end
        if (PRED15_24_buffer[clk] != PRED15_24_buffer[!clk]) begin
          $fwrite(f, "Register (15,24) Value: %h\n", PRED15_24_buffer[clk]);
        end
        if (PRED15_25_buffer[clk] != PRED15_25_buffer[!clk]) begin
          $fwrite(f, "Register (15,25) Value: %h\n", PRED15_25_buffer[clk]);
        end
        if (PRED15_26_buffer[clk] != PRED15_26_buffer[!clk]) begin
          $fwrite(f, "Register (15,26) Value: %h\n", PRED15_26_buffer[clk]);
        end
        if (PRED15_27_buffer[clk] != PRED15_27_buffer[!clk]) begin
          $fwrite(f, "Register (15,27) Value: %h\n", PRED15_27_buffer[clk]);
        end
        if (PRED15_28_buffer[clk] != PRED15_28_buffer[!clk]) begin
          $fwrite(f, "Register (15,28) Value: %h\n", PRED15_28_buffer[clk]);
        end
        if (PRED15_29_buffer[clk] != PRED15_29_buffer[!clk]) begin
          $fwrite(f, "Register (15,29) Value: %h\n", PRED15_29_buffer[clk]);
        end
        if (PRED15_30_buffer[clk] != PRED15_30_buffer[!clk]) begin
          $fwrite(f, "Register (15,30) Value: %h\n", PRED15_30_buffer[clk]);
        end
        if (PRED15_31_buffer[clk] != PRED15_31_buffer[!clk]) begin
          $fwrite(f, "Register (15,31) Value: %h\n", PRED15_31_buffer[clk]);
        end
        if (PRED16_0_buffer[clk] != PRED16_0_buffer[!clk]) begin
          $fwrite(f, "Register (16,0) Value: %h\n", PRED16_0_buffer[clk]);
        end
        if (PRED16_1_buffer[clk] != PRED16_1_buffer[!clk]) begin
          $fwrite(f, "Register (16,1) Value: %h\n", PRED16_1_buffer[clk]);
        end
        if (PRED16_2_buffer[clk] != PRED16_2_buffer[!clk]) begin
          $fwrite(f, "Register (16,2) Value: %h\n", PRED16_2_buffer[clk]);
        end
        if (PRED16_3_buffer[clk] != PRED16_3_buffer[!clk]) begin
          $fwrite(f, "Register (16,3) Value: %h\n", PRED16_3_buffer[clk]);
        end
        if (PRED16_4_buffer[clk] != PRED16_4_buffer[!clk]) begin
          $fwrite(f, "Register (16,4) Value: %h\n", PRED16_4_buffer[clk]);
        end
        if (PRED16_5_buffer[clk] != PRED16_5_buffer[!clk]) begin
          $fwrite(f, "Register (16,5) Value: %h\n", PRED16_5_buffer[clk]);
        end
        if (PRED16_6_buffer[clk] != PRED16_6_buffer[!clk]) begin
          $fwrite(f, "Register (16,6) Value: %h\n", PRED16_6_buffer[clk]);
        end
        if (PRED16_7_buffer[clk] != PRED16_7_buffer[!clk]) begin
          $fwrite(f, "Register (16,7) Value: %h\n", PRED16_7_buffer[clk]);
        end
        if (PRED16_8_buffer[clk] != PRED16_8_buffer[!clk]) begin
          $fwrite(f, "Register (16,8) Value: %h\n", PRED16_8_buffer[clk]);
        end
        if (PRED16_9_buffer[clk] != PRED16_9_buffer[!clk]) begin
          $fwrite(f, "Register (16,9) Value: %h\n", PRED16_9_buffer[clk]);
        end
        if (PRED16_10_buffer[clk] != PRED16_10_buffer[!clk]) begin
          $fwrite(f, "Register (16,10) Value: %h\n", PRED16_10_buffer[clk]);
        end
        if (PRED16_11_buffer[clk] != PRED16_11_buffer[!clk]) begin
          $fwrite(f, "Register (16,11) Value: %h\n", PRED16_11_buffer[clk]);
        end
        if (PRED16_12_buffer[clk] != PRED16_12_buffer[!clk]) begin
          $fwrite(f, "Register (16,12) Value: %h\n", PRED16_12_buffer[clk]);
        end
        if (PRED16_13_buffer[clk] != PRED16_13_buffer[!clk]) begin
          $fwrite(f, "Register (16,13) Value: %h\n", PRED16_13_buffer[clk]);
        end
        if (PRED16_14_buffer[clk] != PRED16_14_buffer[!clk]) begin
          $fwrite(f, "Register (16,14) Value: %h\n", PRED16_14_buffer[clk]);
        end
        if (PRED16_15_buffer[clk] != PRED16_15_buffer[!clk]) begin
          $fwrite(f, "Register (16,15) Value: %h\n", PRED16_15_buffer[clk]);
        end
        if (PRED16_16_buffer[clk] != PRED16_16_buffer[!clk]) begin
          $fwrite(f, "Register (16,16) Value: %h\n", PRED16_16_buffer[clk]);
        end
        if (PRED16_17_buffer[clk] != PRED16_17_buffer[!clk]) begin
          $fwrite(f, "Register (16,17) Value: %h\n", PRED16_17_buffer[clk]);
        end
        if (PRED16_18_buffer[clk] != PRED16_18_buffer[!clk]) begin
          $fwrite(f, "Register (16,18) Value: %h\n", PRED16_18_buffer[clk]);
        end
        if (PRED16_19_buffer[clk] != PRED16_19_buffer[!clk]) begin
          $fwrite(f, "Register (16,19) Value: %h\n", PRED16_19_buffer[clk]);
        end
        if (PRED16_20_buffer[clk] != PRED16_20_buffer[!clk]) begin
          $fwrite(f, "Register (16,20) Value: %h\n", PRED16_20_buffer[clk]);
        end
        if (PRED16_21_buffer[clk] != PRED16_21_buffer[!clk]) begin
          $fwrite(f, "Register (16,21) Value: %h\n", PRED16_21_buffer[clk]);
        end
        if (PRED16_22_buffer[clk] != PRED16_22_buffer[!clk]) begin
          $fwrite(f, "Register (16,22) Value: %h\n", PRED16_22_buffer[clk]);
        end
        if (PRED16_23_buffer[clk] != PRED16_23_buffer[!clk]) begin
          $fwrite(f, "Register (16,23) Value: %h\n", PRED16_23_buffer[clk]);
        end
        if (PRED16_24_buffer[clk] != PRED16_24_buffer[!clk]) begin
          $fwrite(f, "Register (16,24) Value: %h\n", PRED16_24_buffer[clk]);
        end
        if (PRED16_25_buffer[clk] != PRED16_25_buffer[!clk]) begin
          $fwrite(f, "Register (16,25) Value: %h\n", PRED16_25_buffer[clk]);
        end
        if (PRED16_26_buffer[clk] != PRED16_26_buffer[!clk]) begin
          $fwrite(f, "Register (16,26) Value: %h\n", PRED16_26_buffer[clk]);
        end
        if (PRED16_27_buffer[clk] != PRED16_27_buffer[!clk]) begin
          $fwrite(f, "Register (16,27) Value: %h\n", PRED16_27_buffer[clk]);
        end
        if (PRED16_28_buffer[clk] != PRED16_28_buffer[!clk]) begin
          $fwrite(f, "Register (16,28) Value: %h\n", PRED16_28_buffer[clk]);
        end
        if (PRED16_29_buffer[clk] != PRED16_29_buffer[!clk]) begin
          $fwrite(f, "Register (16,29) Value: %h\n", PRED16_29_buffer[clk]);
        end
        if (PRED16_30_buffer[clk] != PRED16_30_buffer[!clk]) begin
          $fwrite(f, "Register (16,30) Value: %h\n", PRED16_30_buffer[clk]);
        end
        if (PRED16_31_buffer[clk] != PRED16_31_buffer[!clk]) begin
          $fwrite(f, "Register (16,31) Value: %h\n", PRED16_31_buffer[clk]);
        end
        if (PRED17_0_buffer[clk] != PRED17_0_buffer[!clk]) begin
          $fwrite(f, "Register (17,0) Value: %h\n", PRED17_0_buffer[clk]);
        end
        if (PRED17_1_buffer[clk] != PRED17_1_buffer[!clk]) begin
          $fwrite(f, "Register (17,1) Value: %h\n", PRED17_1_buffer[clk]);
        end
        if (PRED17_2_buffer[clk] != PRED17_2_buffer[!clk]) begin
          $fwrite(f, "Register (17,2) Value: %h\n", PRED17_2_buffer[clk]);
        end
        if (PRED17_3_buffer[clk] != PRED17_3_buffer[!clk]) begin
          $fwrite(f, "Register (17,3) Value: %h\n", PRED17_3_buffer[clk]);
        end
        if (PRED17_4_buffer[clk] != PRED17_4_buffer[!clk]) begin
          $fwrite(f, "Register (17,4) Value: %h\n", PRED17_4_buffer[clk]);
        end
        if (PRED17_5_buffer[clk] != PRED17_5_buffer[!clk]) begin
          $fwrite(f, "Register (17,5) Value: %h\n", PRED17_5_buffer[clk]);
        end
        if (PRED17_6_buffer[clk] != PRED17_6_buffer[!clk]) begin
          $fwrite(f, "Register (17,6) Value: %h\n", PRED17_6_buffer[clk]);
        end
        if (PRED17_7_buffer[clk] != PRED17_7_buffer[!clk]) begin
          $fwrite(f, "Register (17,7) Value: %h\n", PRED17_7_buffer[clk]);
        end
        if (PRED17_8_buffer[clk] != PRED17_8_buffer[!clk]) begin
          $fwrite(f, "Register (17,8) Value: %h\n", PRED17_8_buffer[clk]);
        end
        if (PRED17_9_buffer[clk] != PRED17_9_buffer[!clk]) begin
          $fwrite(f, "Register (17,9) Value: %h\n", PRED17_9_buffer[clk]);
        end
        if (PRED17_10_buffer[clk] != PRED17_10_buffer[!clk]) begin
          $fwrite(f, "Register (17,10) Value: %h\n", PRED17_10_buffer[clk]);
        end
        if (PRED17_11_buffer[clk] != PRED17_11_buffer[!clk]) begin
          $fwrite(f, "Register (17,11) Value: %h\n", PRED17_11_buffer[clk]);
        end
        if (PRED17_12_buffer[clk] != PRED17_12_buffer[!clk]) begin
          $fwrite(f, "Register (17,12) Value: %h\n", PRED17_12_buffer[clk]);
        end
        if (PRED17_13_buffer[clk] != PRED17_13_buffer[!clk]) begin
          $fwrite(f, "Register (17,13) Value: %h\n", PRED17_13_buffer[clk]);
        end
        if (PRED17_14_buffer[clk] != PRED17_14_buffer[!clk]) begin
          $fwrite(f, "Register (17,14) Value: %h\n", PRED17_14_buffer[clk]);
        end
        if (PRED17_15_buffer[clk] != PRED17_15_buffer[!clk]) begin
          $fwrite(f, "Register (17,15) Value: %h\n", PRED17_15_buffer[clk]);
        end
        if (PRED17_16_buffer[clk] != PRED17_16_buffer[!clk]) begin
          $fwrite(f, "Register (17,16) Value: %h\n", PRED17_16_buffer[clk]);
        end
        if (PRED17_17_buffer[clk] != PRED17_17_buffer[!clk]) begin
          $fwrite(f, "Register (17,17) Value: %h\n", PRED17_17_buffer[clk]);
        end
        if (PRED17_18_buffer[clk] != PRED17_18_buffer[!clk]) begin
          $fwrite(f, "Register (17,18) Value: %h\n", PRED17_18_buffer[clk]);
        end
        if (PRED17_19_buffer[clk] != PRED17_19_buffer[!clk]) begin
          $fwrite(f, "Register (17,19) Value: %h\n", PRED17_19_buffer[clk]);
        end
        if (PRED17_20_buffer[clk] != PRED17_20_buffer[!clk]) begin
          $fwrite(f, "Register (17,20) Value: %h\n", PRED17_20_buffer[clk]);
        end
        if (PRED17_21_buffer[clk] != PRED17_21_buffer[!clk]) begin
          $fwrite(f, "Register (17,21) Value: %h\n", PRED17_21_buffer[clk]);
        end
        if (PRED17_22_buffer[clk] != PRED17_22_buffer[!clk]) begin
          $fwrite(f, "Register (17,22) Value: %h\n", PRED17_22_buffer[clk]);
        end
        if (PRED17_23_buffer[clk] != PRED17_23_buffer[!clk]) begin
          $fwrite(f, "Register (17,23) Value: %h\n", PRED17_23_buffer[clk]);
        end
        if (PRED17_24_buffer[clk] != PRED17_24_buffer[!clk]) begin
          $fwrite(f, "Register (17,24) Value: %h\n", PRED17_24_buffer[clk]);
        end
        if (PRED17_25_buffer[clk] != PRED17_25_buffer[!clk]) begin
          $fwrite(f, "Register (17,25) Value: %h\n", PRED17_25_buffer[clk]);
        end
        if (PRED17_26_buffer[clk] != PRED17_26_buffer[!clk]) begin
          $fwrite(f, "Register (17,26) Value: %h\n", PRED17_26_buffer[clk]);
        end
        if (PRED17_27_buffer[clk] != PRED17_27_buffer[!clk]) begin
          $fwrite(f, "Register (17,27) Value: %h\n", PRED17_27_buffer[clk]);
        end
        if (PRED17_28_buffer[clk] != PRED17_28_buffer[!clk]) begin
          $fwrite(f, "Register (17,28) Value: %h\n", PRED17_28_buffer[clk]);
        end
        if (PRED17_29_buffer[clk] != PRED17_29_buffer[!clk]) begin
          $fwrite(f, "Register (17,29) Value: %h\n", PRED17_29_buffer[clk]);
        end
        if (PRED17_30_buffer[clk] != PRED17_30_buffer[!clk]) begin
          $fwrite(f, "Register (17,30) Value: %h\n", PRED17_30_buffer[clk]);
        end
        if (PRED17_31_buffer[clk] != PRED17_31_buffer[!clk]) begin
          $fwrite(f, "Register (17,31) Value: %h\n", PRED17_31_buffer[clk]);
        end
        if (PRED18_0_buffer[clk] != PRED18_0_buffer[!clk]) begin
          $fwrite(f, "Register (18,0) Value: %h\n", PRED18_0_buffer[clk]);
        end
        if (PRED18_1_buffer[clk] != PRED18_1_buffer[!clk]) begin
          $fwrite(f, "Register (18,1) Value: %h\n", PRED18_1_buffer[clk]);
        end
        if (PRED18_2_buffer[clk] != PRED18_2_buffer[!clk]) begin
          $fwrite(f, "Register (18,2) Value: %h\n", PRED18_2_buffer[clk]);
        end
        if (PRED18_3_buffer[clk] != PRED18_3_buffer[!clk]) begin
          $fwrite(f, "Register (18,3) Value: %h\n", PRED18_3_buffer[clk]);
        end
        if (PRED18_4_buffer[clk] != PRED18_4_buffer[!clk]) begin
          $fwrite(f, "Register (18,4) Value: %h\n", PRED18_4_buffer[clk]);
        end
        if (PRED18_5_buffer[clk] != PRED18_5_buffer[!clk]) begin
          $fwrite(f, "Register (18,5) Value: %h\n", PRED18_5_buffer[clk]);
        end
        if (PRED18_6_buffer[clk] != PRED18_6_buffer[!clk]) begin
          $fwrite(f, "Register (18,6) Value: %h\n", PRED18_6_buffer[clk]);
        end
        if (PRED18_7_buffer[clk] != PRED18_7_buffer[!clk]) begin
          $fwrite(f, "Register (18,7) Value: %h\n", PRED18_7_buffer[clk]);
        end
        if (PRED18_8_buffer[clk] != PRED18_8_buffer[!clk]) begin
          $fwrite(f, "Register (18,8) Value: %h\n", PRED18_8_buffer[clk]);
        end
        if (PRED18_9_buffer[clk] != PRED18_9_buffer[!clk]) begin
          $fwrite(f, "Register (18,9) Value: %h\n", PRED18_9_buffer[clk]);
        end
        if (PRED18_10_buffer[clk] != PRED18_10_buffer[!clk]) begin
          $fwrite(f, "Register (18,10) Value: %h\n", PRED18_10_buffer[clk]);
        end
        if (PRED18_11_buffer[clk] != PRED18_11_buffer[!clk]) begin
          $fwrite(f, "Register (18,11) Value: %h\n", PRED18_11_buffer[clk]);
        end
        if (PRED18_12_buffer[clk] != PRED18_12_buffer[!clk]) begin
          $fwrite(f, "Register (18,12) Value: %h\n", PRED18_12_buffer[clk]);
        end
        if (PRED18_13_buffer[clk] != PRED18_13_buffer[!clk]) begin
          $fwrite(f, "Register (18,13) Value: %h\n", PRED18_13_buffer[clk]);
        end
        if (PRED18_14_buffer[clk] != PRED18_14_buffer[!clk]) begin
          $fwrite(f, "Register (18,14) Value: %h\n", PRED18_14_buffer[clk]);
        end
        if (PRED18_15_buffer[clk] != PRED18_15_buffer[!clk]) begin
          $fwrite(f, "Register (18,15) Value: %h\n", PRED18_15_buffer[clk]);
        end
        if (PRED18_16_buffer[clk] != PRED18_16_buffer[!clk]) begin
          $fwrite(f, "Register (18,16) Value: %h\n", PRED18_16_buffer[clk]);
        end
        if (PRED18_17_buffer[clk] != PRED18_17_buffer[!clk]) begin
          $fwrite(f, "Register (18,17) Value: %h\n", PRED18_17_buffer[clk]);
        end
        if (PRED18_18_buffer[clk] != PRED18_18_buffer[!clk]) begin
          $fwrite(f, "Register (18,18) Value: %h\n", PRED18_18_buffer[clk]);
        end
        if (PRED18_19_buffer[clk] != PRED18_19_buffer[!clk]) begin
          $fwrite(f, "Register (18,19) Value: %h\n", PRED18_19_buffer[clk]);
        end
        if (PRED18_20_buffer[clk] != PRED18_20_buffer[!clk]) begin
          $fwrite(f, "Register (18,20) Value: %h\n", PRED18_20_buffer[clk]);
        end
        if (PRED18_21_buffer[clk] != PRED18_21_buffer[!clk]) begin
          $fwrite(f, "Register (18,21) Value: %h\n", PRED18_21_buffer[clk]);
        end
        if (PRED18_22_buffer[clk] != PRED18_22_buffer[!clk]) begin
          $fwrite(f, "Register (18,22) Value: %h\n", PRED18_22_buffer[clk]);
        end
        if (PRED18_23_buffer[clk] != PRED18_23_buffer[!clk]) begin
          $fwrite(f, "Register (18,23) Value: %h\n", PRED18_23_buffer[clk]);
        end
        if (PRED18_24_buffer[clk] != PRED18_24_buffer[!clk]) begin
          $fwrite(f, "Register (18,24) Value: %h\n", PRED18_24_buffer[clk]);
        end
        if (PRED18_25_buffer[clk] != PRED18_25_buffer[!clk]) begin
          $fwrite(f, "Register (18,25) Value: %h\n", PRED18_25_buffer[clk]);
        end
        if (PRED18_26_buffer[clk] != PRED18_26_buffer[!clk]) begin
          $fwrite(f, "Register (18,26) Value: %h\n", PRED18_26_buffer[clk]);
        end
        if (PRED18_27_buffer[clk] != PRED18_27_buffer[!clk]) begin
          $fwrite(f, "Register (18,27) Value: %h\n", PRED18_27_buffer[clk]);
        end
        if (PRED18_28_buffer[clk] != PRED18_28_buffer[!clk]) begin
          $fwrite(f, "Register (18,28) Value: %h\n", PRED18_28_buffer[clk]);
        end
        if (PRED18_29_buffer[clk] != PRED18_29_buffer[!clk]) begin
          $fwrite(f, "Register (18,29) Value: %h\n", PRED18_29_buffer[clk]);
        end
        if (PRED18_30_buffer[clk] != PRED18_30_buffer[!clk]) begin
          $fwrite(f, "Register (18,30) Value: %h\n", PRED18_30_buffer[clk]);
        end
        if (PRED18_31_buffer[clk] != PRED18_31_buffer[!clk]) begin
          $fwrite(f, "Register (18,31) Value: %h\n", PRED18_31_buffer[clk]);
        end
        if (PRED19_0_buffer[clk] != PRED19_0_buffer[!clk]) begin
          $fwrite(f, "Register (19,0) Value: %h\n", PRED19_0_buffer[clk]);
        end
        if (PRED19_1_buffer[clk] != PRED19_1_buffer[!clk]) begin
          $fwrite(f, "Register (19,1) Value: %h\n", PRED19_1_buffer[clk]);
        end
        if (PRED19_2_buffer[clk] != PRED19_2_buffer[!clk]) begin
          $fwrite(f, "Register (19,2) Value: %h\n", PRED19_2_buffer[clk]);
        end
        if (PRED19_3_buffer[clk] != PRED19_3_buffer[!clk]) begin
          $fwrite(f, "Register (19,3) Value: %h\n", PRED19_3_buffer[clk]);
        end
        if (PRED19_4_buffer[clk] != PRED19_4_buffer[!clk]) begin
          $fwrite(f, "Register (19,4) Value: %h\n", PRED19_4_buffer[clk]);
        end
        if (PRED19_5_buffer[clk] != PRED19_5_buffer[!clk]) begin
          $fwrite(f, "Register (19,5) Value: %h\n", PRED19_5_buffer[clk]);
        end
        if (PRED19_6_buffer[clk] != PRED19_6_buffer[!clk]) begin
          $fwrite(f, "Register (19,6) Value: %h\n", PRED19_6_buffer[clk]);
        end
        if (PRED19_7_buffer[clk] != PRED19_7_buffer[!clk]) begin
          $fwrite(f, "Register (19,7) Value: %h\n", PRED19_7_buffer[clk]);
        end
        if (PRED19_8_buffer[clk] != PRED19_8_buffer[!clk]) begin
          $fwrite(f, "Register (19,8) Value: %h\n", PRED19_8_buffer[clk]);
        end
        if (PRED19_9_buffer[clk] != PRED19_9_buffer[!clk]) begin
          $fwrite(f, "Register (19,9) Value: %h\n", PRED19_9_buffer[clk]);
        end
        if (PRED19_10_buffer[clk] != PRED19_10_buffer[!clk]) begin
          $fwrite(f, "Register (19,10) Value: %h\n", PRED19_10_buffer[clk]);
        end
        if (PRED19_11_buffer[clk] != PRED19_11_buffer[!clk]) begin
          $fwrite(f, "Register (19,11) Value: %h\n", PRED19_11_buffer[clk]);
        end
        if (PRED19_12_buffer[clk] != PRED19_12_buffer[!clk]) begin
          $fwrite(f, "Register (19,12) Value: %h\n", PRED19_12_buffer[clk]);
        end
        if (PRED19_13_buffer[clk] != PRED19_13_buffer[!clk]) begin
          $fwrite(f, "Register (19,13) Value: %h\n", PRED19_13_buffer[clk]);
        end
        if (PRED19_14_buffer[clk] != PRED19_14_buffer[!clk]) begin
          $fwrite(f, "Register (19,14) Value: %h\n", PRED19_14_buffer[clk]);
        end
        if (PRED19_15_buffer[clk] != PRED19_15_buffer[!clk]) begin
          $fwrite(f, "Register (19,15) Value: %h\n", PRED19_15_buffer[clk]);
        end
        if (PRED19_16_buffer[clk] != PRED19_16_buffer[!clk]) begin
          $fwrite(f, "Register (19,16) Value: %h\n", PRED19_16_buffer[clk]);
        end
        if (PRED19_17_buffer[clk] != PRED19_17_buffer[!clk]) begin
          $fwrite(f, "Register (19,17) Value: %h\n", PRED19_17_buffer[clk]);
        end
        if (PRED19_18_buffer[clk] != PRED19_18_buffer[!clk]) begin
          $fwrite(f, "Register (19,18) Value: %h\n", PRED19_18_buffer[clk]);
        end
        if (PRED19_19_buffer[clk] != PRED19_19_buffer[!clk]) begin
          $fwrite(f, "Register (19,19) Value: %h\n", PRED19_19_buffer[clk]);
        end
        if (PRED19_20_buffer[clk] != PRED19_20_buffer[!clk]) begin
          $fwrite(f, "Register (19,20) Value: %h\n", PRED19_20_buffer[clk]);
        end
        if (PRED19_21_buffer[clk] != PRED19_21_buffer[!clk]) begin
          $fwrite(f, "Register (19,21) Value: %h\n", PRED19_21_buffer[clk]);
        end
        if (PRED19_22_buffer[clk] != PRED19_22_buffer[!clk]) begin
          $fwrite(f, "Register (19,22) Value: %h\n", PRED19_22_buffer[clk]);
        end
        if (PRED19_23_buffer[clk] != PRED19_23_buffer[!clk]) begin
          $fwrite(f, "Register (19,23) Value: %h\n", PRED19_23_buffer[clk]);
        end
        if (PRED19_24_buffer[clk] != PRED19_24_buffer[!clk]) begin
          $fwrite(f, "Register (19,24) Value: %h\n", PRED19_24_buffer[clk]);
        end
        if (PRED19_25_buffer[clk] != PRED19_25_buffer[!clk]) begin
          $fwrite(f, "Register (19,25) Value: %h\n", PRED19_25_buffer[clk]);
        end
        if (PRED19_26_buffer[clk] != PRED19_26_buffer[!clk]) begin
          $fwrite(f, "Register (19,26) Value: %h\n", PRED19_26_buffer[clk]);
        end
        if (PRED19_27_buffer[clk] != PRED19_27_buffer[!clk]) begin
          $fwrite(f, "Register (19,27) Value: %h\n", PRED19_27_buffer[clk]);
        end
        if (PRED19_28_buffer[clk] != PRED19_28_buffer[!clk]) begin
          $fwrite(f, "Register (19,28) Value: %h\n", PRED19_28_buffer[clk]);
        end
        if (PRED19_29_buffer[clk] != PRED19_29_buffer[!clk]) begin
          $fwrite(f, "Register (19,29) Value: %h\n", PRED19_29_buffer[clk]);
        end
        if (PRED19_30_buffer[clk] != PRED19_30_buffer[!clk]) begin
          $fwrite(f, "Register (19,30) Value: %h\n", PRED19_30_buffer[clk]);
        end
        if (PRED19_31_buffer[clk] != PRED19_31_buffer[!clk]) begin
          $fwrite(f, "Register (19,31) Value: %h\n", PRED19_31_buffer[clk]);
        end
        if (PRED20_0_buffer[clk] != PRED20_0_buffer[!clk]) begin
          $fwrite(f, "Register (20,0) Value: %h\n", PRED20_0_buffer[clk]);
        end
        if (PRED20_1_buffer[clk] != PRED20_1_buffer[!clk]) begin
          $fwrite(f, "Register (20,1) Value: %h\n", PRED20_1_buffer[clk]);
        end
        if (PRED20_2_buffer[clk] != PRED20_2_buffer[!clk]) begin
          $fwrite(f, "Register (20,2) Value: %h\n", PRED20_2_buffer[clk]);
        end
        if (PRED20_3_buffer[clk] != PRED20_3_buffer[!clk]) begin
          $fwrite(f, "Register (20,3) Value: %h\n", PRED20_3_buffer[clk]);
        end
        if (PRED20_4_buffer[clk] != PRED20_4_buffer[!clk]) begin
          $fwrite(f, "Register (20,4) Value: %h\n", PRED20_4_buffer[clk]);
        end
        if (PRED20_5_buffer[clk] != PRED20_5_buffer[!clk]) begin
          $fwrite(f, "Register (20,5) Value: %h\n", PRED20_5_buffer[clk]);
        end
        if (PRED20_6_buffer[clk] != PRED20_6_buffer[!clk]) begin
          $fwrite(f, "Register (20,6) Value: %h\n", PRED20_6_buffer[clk]);
        end
        if (PRED20_7_buffer[clk] != PRED20_7_buffer[!clk]) begin
          $fwrite(f, "Register (20,7) Value: %h\n", PRED20_7_buffer[clk]);
        end
        if (PRED20_8_buffer[clk] != PRED20_8_buffer[!clk]) begin
          $fwrite(f, "Register (20,8) Value: %h\n", PRED20_8_buffer[clk]);
        end
        if (PRED20_9_buffer[clk] != PRED20_9_buffer[!clk]) begin
          $fwrite(f, "Register (20,9) Value: %h\n", PRED20_9_buffer[clk]);
        end
        if (PRED20_10_buffer[clk] != PRED20_10_buffer[!clk]) begin
          $fwrite(f, "Register (20,10) Value: %h\n", PRED20_10_buffer[clk]);
        end
        if (PRED20_11_buffer[clk] != PRED20_11_buffer[!clk]) begin
          $fwrite(f, "Register (20,11) Value: %h\n", PRED20_11_buffer[clk]);
        end
        if (PRED20_12_buffer[clk] != PRED20_12_buffer[!clk]) begin
          $fwrite(f, "Register (20,12) Value: %h\n", PRED20_12_buffer[clk]);
        end
        if (PRED20_13_buffer[clk] != PRED20_13_buffer[!clk]) begin
          $fwrite(f, "Register (20,13) Value: %h\n", PRED20_13_buffer[clk]);
        end
        if (PRED20_14_buffer[clk] != PRED20_14_buffer[!clk]) begin
          $fwrite(f, "Register (20,14) Value: %h\n", PRED20_14_buffer[clk]);
        end
        if (PRED20_15_buffer[clk] != PRED20_15_buffer[!clk]) begin
          $fwrite(f, "Register (20,15) Value: %h\n", PRED20_15_buffer[clk]);
        end
        if (PRED20_16_buffer[clk] != PRED20_16_buffer[!clk]) begin
          $fwrite(f, "Register (20,16) Value: %h\n", PRED20_16_buffer[clk]);
        end
        if (PRED20_17_buffer[clk] != PRED20_17_buffer[!clk]) begin
          $fwrite(f, "Register (20,17) Value: %h\n", PRED20_17_buffer[clk]);
        end
        if (PRED20_18_buffer[clk] != PRED20_18_buffer[!clk]) begin
          $fwrite(f, "Register (20,18) Value: %h\n", PRED20_18_buffer[clk]);
        end
        if (PRED20_19_buffer[clk] != PRED20_19_buffer[!clk]) begin
          $fwrite(f, "Register (20,19) Value: %h\n", PRED20_19_buffer[clk]);
        end
        if (PRED20_20_buffer[clk] != PRED20_20_buffer[!clk]) begin
          $fwrite(f, "Register (20,20) Value: %h\n", PRED20_20_buffer[clk]);
        end
        if (PRED20_21_buffer[clk] != PRED20_21_buffer[!clk]) begin
          $fwrite(f, "Register (20,21) Value: %h\n", PRED20_21_buffer[clk]);
        end
        if (PRED20_22_buffer[clk] != PRED20_22_buffer[!clk]) begin
          $fwrite(f, "Register (20,22) Value: %h\n", PRED20_22_buffer[clk]);
        end
        if (PRED20_23_buffer[clk] != PRED20_23_buffer[!clk]) begin
          $fwrite(f, "Register (20,23) Value: %h\n", PRED20_23_buffer[clk]);
        end
        if (PRED20_24_buffer[clk] != PRED20_24_buffer[!clk]) begin
          $fwrite(f, "Register (20,24) Value: %h\n", PRED20_24_buffer[clk]);
        end
        if (PRED20_25_buffer[clk] != PRED20_25_buffer[!clk]) begin
          $fwrite(f, "Register (20,25) Value: %h\n", PRED20_25_buffer[clk]);
        end
        if (PRED20_26_buffer[clk] != PRED20_26_buffer[!clk]) begin
          $fwrite(f, "Register (20,26) Value: %h\n", PRED20_26_buffer[clk]);
        end
        if (PRED20_27_buffer[clk] != PRED20_27_buffer[!clk]) begin
          $fwrite(f, "Register (20,27) Value: %h\n", PRED20_27_buffer[clk]);
        end
        if (PRED20_28_buffer[clk] != PRED20_28_buffer[!clk]) begin
          $fwrite(f, "Register (20,28) Value: %h\n", PRED20_28_buffer[clk]);
        end
        if (PRED20_29_buffer[clk] != PRED20_29_buffer[!clk]) begin
          $fwrite(f, "Register (20,29) Value: %h\n", PRED20_29_buffer[clk]);
        end
        if (PRED20_30_buffer[clk] != PRED20_30_buffer[!clk]) begin
          $fwrite(f, "Register (20,30) Value: %h\n", PRED20_30_buffer[clk]);
        end
        if (PRED20_31_buffer[clk] != PRED20_31_buffer[!clk]) begin
          $fwrite(f, "Register (20,31) Value: %h\n", PRED20_31_buffer[clk]);
        end
        if (PRED21_0_buffer[clk] != PRED21_0_buffer[!clk]) begin
          $fwrite(f, "Register (21,0) Value: %h\n", PRED21_0_buffer[clk]);
        end
        if (PRED21_1_buffer[clk] != PRED21_1_buffer[!clk]) begin
          $fwrite(f, "Register (21,1) Value: %h\n", PRED21_1_buffer[clk]);
        end
        if (PRED21_2_buffer[clk] != PRED21_2_buffer[!clk]) begin
          $fwrite(f, "Register (21,2) Value: %h\n", PRED21_2_buffer[clk]);
        end
        if (PRED21_3_buffer[clk] != PRED21_3_buffer[!clk]) begin
          $fwrite(f, "Register (21,3) Value: %h\n", PRED21_3_buffer[clk]);
        end
        if (PRED21_4_buffer[clk] != PRED21_4_buffer[!clk]) begin
          $fwrite(f, "Register (21,4) Value: %h\n", PRED21_4_buffer[clk]);
        end
        if (PRED21_5_buffer[clk] != PRED21_5_buffer[!clk]) begin
          $fwrite(f, "Register (21,5) Value: %h\n", PRED21_5_buffer[clk]);
        end
        if (PRED21_6_buffer[clk] != PRED21_6_buffer[!clk]) begin
          $fwrite(f, "Register (21,6) Value: %h\n", PRED21_6_buffer[clk]);
        end
        if (PRED21_7_buffer[clk] != PRED21_7_buffer[!clk]) begin
          $fwrite(f, "Register (21,7) Value: %h\n", PRED21_7_buffer[clk]);
        end
        if (PRED21_8_buffer[clk] != PRED21_8_buffer[!clk]) begin
          $fwrite(f, "Register (21,8) Value: %h\n", PRED21_8_buffer[clk]);
        end
        if (PRED21_9_buffer[clk] != PRED21_9_buffer[!clk]) begin
          $fwrite(f, "Register (21,9) Value: %h\n", PRED21_9_buffer[clk]);
        end
        if (PRED21_10_buffer[clk] != PRED21_10_buffer[!clk]) begin
          $fwrite(f, "Register (21,10) Value: %h\n", PRED21_10_buffer[clk]);
        end
        if (PRED21_11_buffer[clk] != PRED21_11_buffer[!clk]) begin
          $fwrite(f, "Register (21,11) Value: %h\n", PRED21_11_buffer[clk]);
        end
        if (PRED21_12_buffer[clk] != PRED21_12_buffer[!clk]) begin
          $fwrite(f, "Register (21,12) Value: %h\n", PRED21_12_buffer[clk]);
        end
        if (PRED21_13_buffer[clk] != PRED21_13_buffer[!clk]) begin
          $fwrite(f, "Register (21,13) Value: %h\n", PRED21_13_buffer[clk]);
        end
        if (PRED21_14_buffer[clk] != PRED21_14_buffer[!clk]) begin
          $fwrite(f, "Register (21,14) Value: %h\n", PRED21_14_buffer[clk]);
        end
        if (PRED21_15_buffer[clk] != PRED21_15_buffer[!clk]) begin
          $fwrite(f, "Register (21,15) Value: %h\n", PRED21_15_buffer[clk]);
        end
        if (PRED21_16_buffer[clk] != PRED21_16_buffer[!clk]) begin
          $fwrite(f, "Register (21,16) Value: %h\n", PRED21_16_buffer[clk]);
        end
        if (PRED21_17_buffer[clk] != PRED21_17_buffer[!clk]) begin
          $fwrite(f, "Register (21,17) Value: %h\n", PRED21_17_buffer[clk]);
        end
        if (PRED21_18_buffer[clk] != PRED21_18_buffer[!clk]) begin
          $fwrite(f, "Register (21,18) Value: %h\n", PRED21_18_buffer[clk]);
        end
        if (PRED21_19_buffer[clk] != PRED21_19_buffer[!clk]) begin
          $fwrite(f, "Register (21,19) Value: %h\n", PRED21_19_buffer[clk]);
        end
        if (PRED21_20_buffer[clk] != PRED21_20_buffer[!clk]) begin
          $fwrite(f, "Register (21,20) Value: %h\n", PRED21_20_buffer[clk]);
        end
        if (PRED21_21_buffer[clk] != PRED21_21_buffer[!clk]) begin
          $fwrite(f, "Register (21,21) Value: %h\n", PRED21_21_buffer[clk]);
        end
        if (PRED21_22_buffer[clk] != PRED21_22_buffer[!clk]) begin
          $fwrite(f, "Register (21,22) Value: %h\n", PRED21_22_buffer[clk]);
        end
        if (PRED21_23_buffer[clk] != PRED21_23_buffer[!clk]) begin
          $fwrite(f, "Register (21,23) Value: %h\n", PRED21_23_buffer[clk]);
        end
        if (PRED21_24_buffer[clk] != PRED21_24_buffer[!clk]) begin
          $fwrite(f, "Register (21,24) Value: %h\n", PRED21_24_buffer[clk]);
        end
        if (PRED21_25_buffer[clk] != PRED21_25_buffer[!clk]) begin
          $fwrite(f, "Register (21,25) Value: %h\n", PRED21_25_buffer[clk]);
        end
        if (PRED21_26_buffer[clk] != PRED21_26_buffer[!clk]) begin
          $fwrite(f, "Register (21,26) Value: %h\n", PRED21_26_buffer[clk]);
        end
        if (PRED21_27_buffer[clk] != PRED21_27_buffer[!clk]) begin
          $fwrite(f, "Register (21,27) Value: %h\n", PRED21_27_buffer[clk]);
        end
        if (PRED21_28_buffer[clk] != PRED21_28_buffer[!clk]) begin
          $fwrite(f, "Register (21,28) Value: %h\n", PRED21_28_buffer[clk]);
        end
        if (PRED21_29_buffer[clk] != PRED21_29_buffer[!clk]) begin
          $fwrite(f, "Register (21,29) Value: %h\n", PRED21_29_buffer[clk]);
        end
        if (PRED21_30_buffer[clk] != PRED21_30_buffer[!clk]) begin
          $fwrite(f, "Register (21,30) Value: %h\n", PRED21_30_buffer[clk]);
        end
        if (PRED21_31_buffer[clk] != PRED21_31_buffer[!clk]) begin
          $fwrite(f, "Register (21,31) Value: %h\n", PRED21_31_buffer[clk]);
        end
        if (PRED22_0_buffer[clk] != PRED22_0_buffer[!clk]) begin
          $fwrite(f, "Register (22,0) Value: %h\n", PRED22_0_buffer[clk]);
        end
        if (PRED22_1_buffer[clk] != PRED22_1_buffer[!clk]) begin
          $fwrite(f, "Register (22,1) Value: %h\n", PRED22_1_buffer[clk]);
        end
        if (PRED22_2_buffer[clk] != PRED22_2_buffer[!clk]) begin
          $fwrite(f, "Register (22,2) Value: %h\n", PRED22_2_buffer[clk]);
        end
        if (PRED22_3_buffer[clk] != PRED22_3_buffer[!clk]) begin
          $fwrite(f, "Register (22,3) Value: %h\n", PRED22_3_buffer[clk]);
        end
        if (PRED22_4_buffer[clk] != PRED22_4_buffer[!clk]) begin
          $fwrite(f, "Register (22,4) Value: %h\n", PRED22_4_buffer[clk]);
        end
        if (PRED22_5_buffer[clk] != PRED22_5_buffer[!clk]) begin
          $fwrite(f, "Register (22,5) Value: %h\n", PRED22_5_buffer[clk]);
        end
        if (PRED22_6_buffer[clk] != PRED22_6_buffer[!clk]) begin
          $fwrite(f, "Register (22,6) Value: %h\n", PRED22_6_buffer[clk]);
        end
        if (PRED22_7_buffer[clk] != PRED22_7_buffer[!clk]) begin
          $fwrite(f, "Register (22,7) Value: %h\n", PRED22_7_buffer[clk]);
        end
        if (PRED22_8_buffer[clk] != PRED22_8_buffer[!clk]) begin
          $fwrite(f, "Register (22,8) Value: %h\n", PRED22_8_buffer[clk]);
        end
        if (PRED22_9_buffer[clk] != PRED22_9_buffer[!clk]) begin
          $fwrite(f, "Register (22,9) Value: %h\n", PRED22_9_buffer[clk]);
        end
        if (PRED22_10_buffer[clk] != PRED22_10_buffer[!clk]) begin
          $fwrite(f, "Register (22,10) Value: %h\n", PRED22_10_buffer[clk]);
        end
        if (PRED22_11_buffer[clk] != PRED22_11_buffer[!clk]) begin
          $fwrite(f, "Register (22,11) Value: %h\n", PRED22_11_buffer[clk]);
        end
        if (PRED22_12_buffer[clk] != PRED22_12_buffer[!clk]) begin
          $fwrite(f, "Register (22,12) Value: %h\n", PRED22_12_buffer[clk]);
        end
        if (PRED22_13_buffer[clk] != PRED22_13_buffer[!clk]) begin
          $fwrite(f, "Register (22,13) Value: %h\n", PRED22_13_buffer[clk]);
        end
        if (PRED22_14_buffer[clk] != PRED22_14_buffer[!clk]) begin
          $fwrite(f, "Register (22,14) Value: %h\n", PRED22_14_buffer[clk]);
        end
        if (PRED22_15_buffer[clk] != PRED22_15_buffer[!clk]) begin
          $fwrite(f, "Register (22,15) Value: %h\n", PRED22_15_buffer[clk]);
        end
        if (PRED22_16_buffer[clk] != PRED22_16_buffer[!clk]) begin
          $fwrite(f, "Register (22,16) Value: %h\n", PRED22_16_buffer[clk]);
        end
        if (PRED22_17_buffer[clk] != PRED22_17_buffer[!clk]) begin
          $fwrite(f, "Register (22,17) Value: %h\n", PRED22_17_buffer[clk]);
        end
        if (PRED22_18_buffer[clk] != PRED22_18_buffer[!clk]) begin
          $fwrite(f, "Register (22,18) Value: %h\n", PRED22_18_buffer[clk]);
        end
        if (PRED22_19_buffer[clk] != PRED22_19_buffer[!clk]) begin
          $fwrite(f, "Register (22,19) Value: %h\n", PRED22_19_buffer[clk]);
        end
        if (PRED22_20_buffer[clk] != PRED22_20_buffer[!clk]) begin
          $fwrite(f, "Register (22,20) Value: %h\n", PRED22_20_buffer[clk]);
        end
        if (PRED22_21_buffer[clk] != PRED22_21_buffer[!clk]) begin
          $fwrite(f, "Register (22,21) Value: %h\n", PRED22_21_buffer[clk]);
        end
        if (PRED22_22_buffer[clk] != PRED22_22_buffer[!clk]) begin
          $fwrite(f, "Register (22,22) Value: %h\n", PRED22_22_buffer[clk]);
        end
        if (PRED22_23_buffer[clk] != PRED22_23_buffer[!clk]) begin
          $fwrite(f, "Register (22,23) Value: %h\n", PRED22_23_buffer[clk]);
        end
        if (PRED22_24_buffer[clk] != PRED22_24_buffer[!clk]) begin
          $fwrite(f, "Register (22,24) Value: %h\n", PRED22_24_buffer[clk]);
        end
        if (PRED22_25_buffer[clk] != PRED22_25_buffer[!clk]) begin
          $fwrite(f, "Register (22,25) Value: %h\n", PRED22_25_buffer[clk]);
        end
        if (PRED22_26_buffer[clk] != PRED22_26_buffer[!clk]) begin
          $fwrite(f, "Register (22,26) Value: %h\n", PRED22_26_buffer[clk]);
        end
        if (PRED22_27_buffer[clk] != PRED22_27_buffer[!clk]) begin
          $fwrite(f, "Register (22,27) Value: %h\n", PRED22_27_buffer[clk]);
        end
        if (PRED22_28_buffer[clk] != PRED22_28_buffer[!clk]) begin
          $fwrite(f, "Register (22,28) Value: %h\n", PRED22_28_buffer[clk]);
        end
        if (PRED22_29_buffer[clk] != PRED22_29_buffer[!clk]) begin
          $fwrite(f, "Register (22,29) Value: %h\n", PRED22_29_buffer[clk]);
        end
        if (PRED22_30_buffer[clk] != PRED22_30_buffer[!clk]) begin
          $fwrite(f, "Register (22,30) Value: %h\n", PRED22_30_buffer[clk]);
        end
        if (PRED22_31_buffer[clk] != PRED22_31_buffer[!clk]) begin
          $fwrite(f, "Register (22,31) Value: %h\n", PRED22_31_buffer[clk]);
        end
        if (PRED23_0_buffer[clk] != PRED23_0_buffer[!clk]) begin
          $fwrite(f, "Register (23,0) Value: %h\n", PRED23_0_buffer[clk]);
        end
        if (PRED23_1_buffer[clk] != PRED23_1_buffer[!clk]) begin
          $fwrite(f, "Register (23,1) Value: %h\n", PRED23_1_buffer[clk]);
        end
        if (PRED23_2_buffer[clk] != PRED23_2_buffer[!clk]) begin
          $fwrite(f, "Register (23,2) Value: %h\n", PRED23_2_buffer[clk]);
        end
        if (PRED23_3_buffer[clk] != PRED23_3_buffer[!clk]) begin
          $fwrite(f, "Register (23,3) Value: %h\n", PRED23_3_buffer[clk]);
        end
        if (PRED23_4_buffer[clk] != PRED23_4_buffer[!clk]) begin
          $fwrite(f, "Register (23,4) Value: %h\n", PRED23_4_buffer[clk]);
        end
        if (PRED23_5_buffer[clk] != PRED23_5_buffer[!clk]) begin
          $fwrite(f, "Register (23,5) Value: %h\n", PRED23_5_buffer[clk]);
        end
        if (PRED23_6_buffer[clk] != PRED23_6_buffer[!clk]) begin
          $fwrite(f, "Register (23,6) Value: %h\n", PRED23_6_buffer[clk]);
        end
        if (PRED23_7_buffer[clk] != PRED23_7_buffer[!clk]) begin
          $fwrite(f, "Register (23,7) Value: %h\n", PRED23_7_buffer[clk]);
        end
        if (PRED23_8_buffer[clk] != PRED23_8_buffer[!clk]) begin
          $fwrite(f, "Register (23,8) Value: %h\n", PRED23_8_buffer[clk]);
        end
        if (PRED23_9_buffer[clk] != PRED23_9_buffer[!clk]) begin
          $fwrite(f, "Register (23,9) Value: %h\n", PRED23_9_buffer[clk]);
        end
        if (PRED23_10_buffer[clk] != PRED23_10_buffer[!clk]) begin
          $fwrite(f, "Register (23,10) Value: %h\n", PRED23_10_buffer[clk]);
        end
        if (PRED23_11_buffer[clk] != PRED23_11_buffer[!clk]) begin
          $fwrite(f, "Register (23,11) Value: %h\n", PRED23_11_buffer[clk]);
        end
        if (PRED23_12_buffer[clk] != PRED23_12_buffer[!clk]) begin
          $fwrite(f, "Register (23,12) Value: %h\n", PRED23_12_buffer[clk]);
        end
        if (PRED23_13_buffer[clk] != PRED23_13_buffer[!clk]) begin
          $fwrite(f, "Register (23,13) Value: %h\n", PRED23_13_buffer[clk]);
        end
        if (PRED23_14_buffer[clk] != PRED23_14_buffer[!clk]) begin
          $fwrite(f, "Register (23,14) Value: %h\n", PRED23_14_buffer[clk]);
        end
        if (PRED23_15_buffer[clk] != PRED23_15_buffer[!clk]) begin
          $fwrite(f, "Register (23,15) Value: %h\n", PRED23_15_buffer[clk]);
        end
        if (PRED23_16_buffer[clk] != PRED23_16_buffer[!clk]) begin
          $fwrite(f, "Register (23,16) Value: %h\n", PRED23_16_buffer[clk]);
        end
        if (PRED23_17_buffer[clk] != PRED23_17_buffer[!clk]) begin
          $fwrite(f, "Register (23,17) Value: %h\n", PRED23_17_buffer[clk]);
        end
        if (PRED23_18_buffer[clk] != PRED23_18_buffer[!clk]) begin
          $fwrite(f, "Register (23,18) Value: %h\n", PRED23_18_buffer[clk]);
        end
        if (PRED23_19_buffer[clk] != PRED23_19_buffer[!clk]) begin
          $fwrite(f, "Register (23,19) Value: %h\n", PRED23_19_buffer[clk]);
        end
        if (PRED23_20_buffer[clk] != PRED23_20_buffer[!clk]) begin
          $fwrite(f, "Register (23,20) Value: %h\n", PRED23_20_buffer[clk]);
        end
        if (PRED23_21_buffer[clk] != PRED23_21_buffer[!clk]) begin
          $fwrite(f, "Register (23,21) Value: %h\n", PRED23_21_buffer[clk]);
        end
        if (PRED23_22_buffer[clk] != PRED23_22_buffer[!clk]) begin
          $fwrite(f, "Register (23,22) Value: %h\n", PRED23_22_buffer[clk]);
        end
        if (PRED23_23_buffer[clk] != PRED23_23_buffer[!clk]) begin
          $fwrite(f, "Register (23,23) Value: %h\n", PRED23_23_buffer[clk]);
        end
        if (PRED23_24_buffer[clk] != PRED23_24_buffer[!clk]) begin
          $fwrite(f, "Register (23,24) Value: %h\n", PRED23_24_buffer[clk]);
        end
        if (PRED23_25_buffer[clk] != PRED23_25_buffer[!clk]) begin
          $fwrite(f, "Register (23,25) Value: %h\n", PRED23_25_buffer[clk]);
        end
        if (PRED23_26_buffer[clk] != PRED23_26_buffer[!clk]) begin
          $fwrite(f, "Register (23,26) Value: %h\n", PRED23_26_buffer[clk]);
        end
        if (PRED23_27_buffer[clk] != PRED23_27_buffer[!clk]) begin
          $fwrite(f, "Register (23,27) Value: %h\n", PRED23_27_buffer[clk]);
        end
        if (PRED23_28_buffer[clk] != PRED23_28_buffer[!clk]) begin
          $fwrite(f, "Register (23,28) Value: %h\n", PRED23_28_buffer[clk]);
        end
        if (PRED23_29_buffer[clk] != PRED23_29_buffer[!clk]) begin
          $fwrite(f, "Register (23,29) Value: %h\n", PRED23_29_buffer[clk]);
        end
        if (PRED23_30_buffer[clk] != PRED23_30_buffer[!clk]) begin
          $fwrite(f, "Register (23,30) Value: %h\n", PRED23_30_buffer[clk]);
        end
        if (PRED23_31_buffer[clk] != PRED23_31_buffer[!clk]) begin
          $fwrite(f, "Register (23,31) Value: %h\n", PRED23_31_buffer[clk]);
        end
        if (PRED24_0_buffer[clk] != PRED24_0_buffer[!clk]) begin
          $fwrite(f, "Register (24,0) Value: %h\n", PRED24_0_buffer[clk]);
        end
        if (PRED24_1_buffer[clk] != PRED24_1_buffer[!clk]) begin
          $fwrite(f, "Register (24,1) Value: %h\n", PRED24_1_buffer[clk]);
        end
        if (PRED24_2_buffer[clk] != PRED24_2_buffer[!clk]) begin
          $fwrite(f, "Register (24,2) Value: %h\n", PRED24_2_buffer[clk]);
        end
        if (PRED24_3_buffer[clk] != PRED24_3_buffer[!clk]) begin
          $fwrite(f, "Register (24,3) Value: %h\n", PRED24_3_buffer[clk]);
        end
        if (PRED24_4_buffer[clk] != PRED24_4_buffer[!clk]) begin
          $fwrite(f, "Register (24,4) Value: %h\n", PRED24_4_buffer[clk]);
        end
        if (PRED24_5_buffer[clk] != PRED24_5_buffer[!clk]) begin
          $fwrite(f, "Register (24,5) Value: %h\n", PRED24_5_buffer[clk]);
        end
        if (PRED24_6_buffer[clk] != PRED24_6_buffer[!clk]) begin
          $fwrite(f, "Register (24,6) Value: %h\n", PRED24_6_buffer[clk]);
        end
        if (PRED24_7_buffer[clk] != PRED24_7_buffer[!clk]) begin
          $fwrite(f, "Register (24,7) Value: %h\n", PRED24_7_buffer[clk]);
        end
        if (PRED24_8_buffer[clk] != PRED24_8_buffer[!clk]) begin
          $fwrite(f, "Register (24,8) Value: %h\n", PRED24_8_buffer[clk]);
        end
        if (PRED24_9_buffer[clk] != PRED24_9_buffer[!clk]) begin
          $fwrite(f, "Register (24,9) Value: %h\n", PRED24_9_buffer[clk]);
        end
        if (PRED24_10_buffer[clk] != PRED24_10_buffer[!clk]) begin
          $fwrite(f, "Register (24,10) Value: %h\n", PRED24_10_buffer[clk]);
        end
        if (PRED24_11_buffer[clk] != PRED24_11_buffer[!clk]) begin
          $fwrite(f, "Register (24,11) Value: %h\n", PRED24_11_buffer[clk]);
        end
        if (PRED24_12_buffer[clk] != PRED24_12_buffer[!clk]) begin
          $fwrite(f, "Register (24,12) Value: %h\n", PRED24_12_buffer[clk]);
        end
        if (PRED24_13_buffer[clk] != PRED24_13_buffer[!clk]) begin
          $fwrite(f, "Register (24,13) Value: %h\n", PRED24_13_buffer[clk]);
        end
        if (PRED24_14_buffer[clk] != PRED24_14_buffer[!clk]) begin
          $fwrite(f, "Register (24,14) Value: %h\n", PRED24_14_buffer[clk]);
        end
        if (PRED24_15_buffer[clk] != PRED24_15_buffer[!clk]) begin
          $fwrite(f, "Register (24,15) Value: %h\n", PRED24_15_buffer[clk]);
        end
        if (PRED24_16_buffer[clk] != PRED24_16_buffer[!clk]) begin
          $fwrite(f, "Register (24,16) Value: %h\n", PRED24_16_buffer[clk]);
        end
        if (PRED24_17_buffer[clk] != PRED24_17_buffer[!clk]) begin
          $fwrite(f, "Register (24,17) Value: %h\n", PRED24_17_buffer[clk]);
        end
        if (PRED24_18_buffer[clk] != PRED24_18_buffer[!clk]) begin
          $fwrite(f, "Register (24,18) Value: %h\n", PRED24_18_buffer[clk]);
        end
        if (PRED24_19_buffer[clk] != PRED24_19_buffer[!clk]) begin
          $fwrite(f, "Register (24,19) Value: %h\n", PRED24_19_buffer[clk]);
        end
        if (PRED24_20_buffer[clk] != PRED24_20_buffer[!clk]) begin
          $fwrite(f, "Register (24,20) Value: %h\n", PRED24_20_buffer[clk]);
        end
        if (PRED24_21_buffer[clk] != PRED24_21_buffer[!clk]) begin
          $fwrite(f, "Register (24,21) Value: %h\n", PRED24_21_buffer[clk]);
        end
        if (PRED24_22_buffer[clk] != PRED24_22_buffer[!clk]) begin
          $fwrite(f, "Register (24,22) Value: %h\n", PRED24_22_buffer[clk]);
        end
        if (PRED24_23_buffer[clk] != PRED24_23_buffer[!clk]) begin
          $fwrite(f, "Register (24,23) Value: %h\n", PRED24_23_buffer[clk]);
        end
        if (PRED24_24_buffer[clk] != PRED24_24_buffer[!clk]) begin
          $fwrite(f, "Register (24,24) Value: %h\n", PRED24_24_buffer[clk]);
        end
        if (PRED24_25_buffer[clk] != PRED24_25_buffer[!clk]) begin
          $fwrite(f, "Register (24,25) Value: %h\n", PRED24_25_buffer[clk]);
        end
        if (PRED24_26_buffer[clk] != PRED24_26_buffer[!clk]) begin
          $fwrite(f, "Register (24,26) Value: %h\n", PRED24_26_buffer[clk]);
        end
        if (PRED24_27_buffer[clk] != PRED24_27_buffer[!clk]) begin
          $fwrite(f, "Register (24,27) Value: %h\n", PRED24_27_buffer[clk]);
        end
        if (PRED24_28_buffer[clk] != PRED24_28_buffer[!clk]) begin
          $fwrite(f, "Register (24,28) Value: %h\n", PRED24_28_buffer[clk]);
        end
        if (PRED24_29_buffer[clk] != PRED24_29_buffer[!clk]) begin
          $fwrite(f, "Register (24,29) Value: %h\n", PRED24_29_buffer[clk]);
        end
        if (PRED24_30_buffer[clk] != PRED24_30_buffer[!clk]) begin
          $fwrite(f, "Register (24,30) Value: %h\n", PRED24_30_buffer[clk]);
        end
        if (PRED24_31_buffer[clk] != PRED24_31_buffer[!clk]) begin
          $fwrite(f, "Register (24,31) Value: %h\n", PRED24_31_buffer[clk]);
        end
        if (PRED25_0_buffer[clk] != PRED25_0_buffer[!clk]) begin
          $fwrite(f, "Register (25,0) Value: %h\n", PRED25_0_buffer[clk]);
        end
        if (PRED25_1_buffer[clk] != PRED25_1_buffer[!clk]) begin
          $fwrite(f, "Register (25,1) Value: %h\n", PRED25_1_buffer[clk]);
        end
        if (PRED25_2_buffer[clk] != PRED25_2_buffer[!clk]) begin
          $fwrite(f, "Register (25,2) Value: %h\n", PRED25_2_buffer[clk]);
        end
        if (PRED25_3_buffer[clk] != PRED25_3_buffer[!clk]) begin
          $fwrite(f, "Register (25,3) Value: %h\n", PRED25_3_buffer[clk]);
        end
        if (PRED25_4_buffer[clk] != PRED25_4_buffer[!clk]) begin
          $fwrite(f, "Register (25,4) Value: %h\n", PRED25_4_buffer[clk]);
        end
        if (PRED25_5_buffer[clk] != PRED25_5_buffer[!clk]) begin
          $fwrite(f, "Register (25,5) Value: %h\n", PRED25_5_buffer[clk]);
        end
        if (PRED25_6_buffer[clk] != PRED25_6_buffer[!clk]) begin
          $fwrite(f, "Register (25,6) Value: %h\n", PRED25_6_buffer[clk]);
        end
        if (PRED25_7_buffer[clk] != PRED25_7_buffer[!clk]) begin
          $fwrite(f, "Register (25,7) Value: %h\n", PRED25_7_buffer[clk]);
        end
        if (PRED25_8_buffer[clk] != PRED25_8_buffer[!clk]) begin
          $fwrite(f, "Register (25,8) Value: %h\n", PRED25_8_buffer[clk]);
        end
        if (PRED25_9_buffer[clk] != PRED25_9_buffer[!clk]) begin
          $fwrite(f, "Register (25,9) Value: %h\n", PRED25_9_buffer[clk]);
        end
        if (PRED25_10_buffer[clk] != PRED25_10_buffer[!clk]) begin
          $fwrite(f, "Register (25,10) Value: %h\n", PRED25_10_buffer[clk]);
        end
        if (PRED25_11_buffer[clk] != PRED25_11_buffer[!clk]) begin
          $fwrite(f, "Register (25,11) Value: %h\n", PRED25_11_buffer[clk]);
        end
        if (PRED25_12_buffer[clk] != PRED25_12_buffer[!clk]) begin
          $fwrite(f, "Register (25,12) Value: %h\n", PRED25_12_buffer[clk]);
        end
        if (PRED25_13_buffer[clk] != PRED25_13_buffer[!clk]) begin
          $fwrite(f, "Register (25,13) Value: %h\n", PRED25_13_buffer[clk]);
        end
        if (PRED25_14_buffer[clk] != PRED25_14_buffer[!clk]) begin
          $fwrite(f, "Register (25,14) Value: %h\n", PRED25_14_buffer[clk]);
        end
        if (PRED25_15_buffer[clk] != PRED25_15_buffer[!clk]) begin
          $fwrite(f, "Register (25,15) Value: %h\n", PRED25_15_buffer[clk]);
        end
        if (PRED25_16_buffer[clk] != PRED25_16_buffer[!clk]) begin
          $fwrite(f, "Register (25,16) Value: %h\n", PRED25_16_buffer[clk]);
        end
        if (PRED25_17_buffer[clk] != PRED25_17_buffer[!clk]) begin
          $fwrite(f, "Register (25,17) Value: %h\n", PRED25_17_buffer[clk]);
        end
        if (PRED25_18_buffer[clk] != PRED25_18_buffer[!clk]) begin
          $fwrite(f, "Register (25,18) Value: %h\n", PRED25_18_buffer[clk]);
        end
        if (PRED25_19_buffer[clk] != PRED25_19_buffer[!clk]) begin
          $fwrite(f, "Register (25,19) Value: %h\n", PRED25_19_buffer[clk]);
        end
        if (PRED25_20_buffer[clk] != PRED25_20_buffer[!clk]) begin
          $fwrite(f, "Register (25,20) Value: %h\n", PRED25_20_buffer[clk]);
        end
        if (PRED25_21_buffer[clk] != PRED25_21_buffer[!clk]) begin
          $fwrite(f, "Register (25,21) Value: %h\n", PRED25_21_buffer[clk]);
        end
        if (PRED25_22_buffer[clk] != PRED25_22_buffer[!clk]) begin
          $fwrite(f, "Register (25,22) Value: %h\n", PRED25_22_buffer[clk]);
        end
        if (PRED25_23_buffer[clk] != PRED25_23_buffer[!clk]) begin
          $fwrite(f, "Register (25,23) Value: %h\n", PRED25_23_buffer[clk]);
        end
        if (PRED25_24_buffer[clk] != PRED25_24_buffer[!clk]) begin
          $fwrite(f, "Register (25,24) Value: %h\n", PRED25_24_buffer[clk]);
        end
        if (PRED25_25_buffer[clk] != PRED25_25_buffer[!clk]) begin
          $fwrite(f, "Register (25,25) Value: %h\n", PRED25_25_buffer[clk]);
        end
        if (PRED25_26_buffer[clk] != PRED25_26_buffer[!clk]) begin
          $fwrite(f, "Register (25,26) Value: %h\n", PRED25_26_buffer[clk]);
        end
        if (PRED25_27_buffer[clk] != PRED25_27_buffer[!clk]) begin
          $fwrite(f, "Register (25,27) Value: %h\n", PRED25_27_buffer[clk]);
        end
        if (PRED25_28_buffer[clk] != PRED25_28_buffer[!clk]) begin
          $fwrite(f, "Register (25,28) Value: %h\n", PRED25_28_buffer[clk]);
        end
        if (PRED25_29_buffer[clk] != PRED25_29_buffer[!clk]) begin
          $fwrite(f, "Register (25,29) Value: %h\n", PRED25_29_buffer[clk]);
        end
        if (PRED25_30_buffer[clk] != PRED25_30_buffer[!clk]) begin
          $fwrite(f, "Register (25,30) Value: %h\n", PRED25_30_buffer[clk]);
        end
        if (PRED25_31_buffer[clk] != PRED25_31_buffer[!clk]) begin
          $fwrite(f, "Register (25,31) Value: %h\n", PRED25_31_buffer[clk]);
        end
        if (PRED26_0_buffer[clk] != PRED26_0_buffer[!clk]) begin
          $fwrite(f, "Register (26,0) Value: %h\n", PRED26_0_buffer[clk]);
        end
        if (PRED26_1_buffer[clk] != PRED26_1_buffer[!clk]) begin
          $fwrite(f, "Register (26,1) Value: %h\n", PRED26_1_buffer[clk]);
        end
        if (PRED26_2_buffer[clk] != PRED26_2_buffer[!clk]) begin
          $fwrite(f, "Register (26,2) Value: %h\n", PRED26_2_buffer[clk]);
        end
        if (PRED26_3_buffer[clk] != PRED26_3_buffer[!clk]) begin
          $fwrite(f, "Register (26,3) Value: %h\n", PRED26_3_buffer[clk]);
        end
        if (PRED26_4_buffer[clk] != PRED26_4_buffer[!clk]) begin
          $fwrite(f, "Register (26,4) Value: %h\n", PRED26_4_buffer[clk]);
        end
        if (PRED26_5_buffer[clk] != PRED26_5_buffer[!clk]) begin
          $fwrite(f, "Register (26,5) Value: %h\n", PRED26_5_buffer[clk]);
        end
        if (PRED26_6_buffer[clk] != PRED26_6_buffer[!clk]) begin
          $fwrite(f, "Register (26,6) Value: %h\n", PRED26_6_buffer[clk]);
        end
        if (PRED26_7_buffer[clk] != PRED26_7_buffer[!clk]) begin
          $fwrite(f, "Register (26,7) Value: %h\n", PRED26_7_buffer[clk]);
        end
        if (PRED26_8_buffer[clk] != PRED26_8_buffer[!clk]) begin
          $fwrite(f, "Register (26,8) Value: %h\n", PRED26_8_buffer[clk]);
        end
        if (PRED26_9_buffer[clk] != PRED26_9_buffer[!clk]) begin
          $fwrite(f, "Register (26,9) Value: %h\n", PRED26_9_buffer[clk]);
        end
        if (PRED26_10_buffer[clk] != PRED26_10_buffer[!clk]) begin
          $fwrite(f, "Register (26,10) Value: %h\n", PRED26_10_buffer[clk]);
        end
        if (PRED26_11_buffer[clk] != PRED26_11_buffer[!clk]) begin
          $fwrite(f, "Register (26,11) Value: %h\n", PRED26_11_buffer[clk]);
        end
        if (PRED26_12_buffer[clk] != PRED26_12_buffer[!clk]) begin
          $fwrite(f, "Register (26,12) Value: %h\n", PRED26_12_buffer[clk]);
        end
        if (PRED26_13_buffer[clk] != PRED26_13_buffer[!clk]) begin
          $fwrite(f, "Register (26,13) Value: %h\n", PRED26_13_buffer[clk]);
        end
        if (PRED26_14_buffer[clk] != PRED26_14_buffer[!clk]) begin
          $fwrite(f, "Register (26,14) Value: %h\n", PRED26_14_buffer[clk]);
        end
        if (PRED26_15_buffer[clk] != PRED26_15_buffer[!clk]) begin
          $fwrite(f, "Register (26,15) Value: %h\n", PRED26_15_buffer[clk]);
        end
        if (PRED26_16_buffer[clk] != PRED26_16_buffer[!clk]) begin
          $fwrite(f, "Register (26,16) Value: %h\n", PRED26_16_buffer[clk]);
        end
        if (PRED26_17_buffer[clk] != PRED26_17_buffer[!clk]) begin
          $fwrite(f, "Register (26,17) Value: %h\n", PRED26_17_buffer[clk]);
        end
        if (PRED26_18_buffer[clk] != PRED26_18_buffer[!clk]) begin
          $fwrite(f, "Register (26,18) Value: %h\n", PRED26_18_buffer[clk]);
        end
        if (PRED26_19_buffer[clk] != PRED26_19_buffer[!clk]) begin
          $fwrite(f, "Register (26,19) Value: %h\n", PRED26_19_buffer[clk]);
        end
        if (PRED26_20_buffer[clk] != PRED26_20_buffer[!clk]) begin
          $fwrite(f, "Register (26,20) Value: %h\n", PRED26_20_buffer[clk]);
        end
        if (PRED26_21_buffer[clk] != PRED26_21_buffer[!clk]) begin
          $fwrite(f, "Register (26,21) Value: %h\n", PRED26_21_buffer[clk]);
        end
        if (PRED26_22_buffer[clk] != PRED26_22_buffer[!clk]) begin
          $fwrite(f, "Register (26,22) Value: %h\n", PRED26_22_buffer[clk]);
        end
        if (PRED26_23_buffer[clk] != PRED26_23_buffer[!clk]) begin
          $fwrite(f, "Register (26,23) Value: %h\n", PRED26_23_buffer[clk]);
        end
        if (PRED26_24_buffer[clk] != PRED26_24_buffer[!clk]) begin
          $fwrite(f, "Register (26,24) Value: %h\n", PRED26_24_buffer[clk]);
        end
        if (PRED26_25_buffer[clk] != PRED26_25_buffer[!clk]) begin
          $fwrite(f, "Register (26,25) Value: %h\n", PRED26_25_buffer[clk]);
        end
        if (PRED26_26_buffer[clk] != PRED26_26_buffer[!clk]) begin
          $fwrite(f, "Register (26,26) Value: %h\n", PRED26_26_buffer[clk]);
        end
        if (PRED26_27_buffer[clk] != PRED26_27_buffer[!clk]) begin
          $fwrite(f, "Register (26,27) Value: %h\n", PRED26_27_buffer[clk]);
        end
        if (PRED26_28_buffer[clk] != PRED26_28_buffer[!clk]) begin
          $fwrite(f, "Register (26,28) Value: %h\n", PRED26_28_buffer[clk]);
        end
        if (PRED26_29_buffer[clk] != PRED26_29_buffer[!clk]) begin
          $fwrite(f, "Register (26,29) Value: %h\n", PRED26_29_buffer[clk]);
        end
        if (PRED26_30_buffer[clk] != PRED26_30_buffer[!clk]) begin
          $fwrite(f, "Register (26,30) Value: %h\n", PRED26_30_buffer[clk]);
        end
        if (PRED26_31_buffer[clk] != PRED26_31_buffer[!clk]) begin
          $fwrite(f, "Register (26,31) Value: %h\n", PRED26_31_buffer[clk]);
        end
        if (PRED27_0_buffer[clk] != PRED27_0_buffer[!clk]) begin
          $fwrite(f, "Register (27,0) Value: %h\n", PRED27_0_buffer[clk]);
        end
        if (PRED27_1_buffer[clk] != PRED27_1_buffer[!clk]) begin
          $fwrite(f, "Register (27,1) Value: %h\n", PRED27_1_buffer[clk]);
        end
        if (PRED27_2_buffer[clk] != PRED27_2_buffer[!clk]) begin
          $fwrite(f, "Register (27,2) Value: %h\n", PRED27_2_buffer[clk]);
        end
        if (PRED27_3_buffer[clk] != PRED27_3_buffer[!clk]) begin
          $fwrite(f, "Register (27,3) Value: %h\n", PRED27_3_buffer[clk]);
        end
        if (PRED27_4_buffer[clk] != PRED27_4_buffer[!clk]) begin
          $fwrite(f, "Register (27,4) Value: %h\n", PRED27_4_buffer[clk]);
        end
        if (PRED27_5_buffer[clk] != PRED27_5_buffer[!clk]) begin
          $fwrite(f, "Register (27,5) Value: %h\n", PRED27_5_buffer[clk]);
        end
        if (PRED27_6_buffer[clk] != PRED27_6_buffer[!clk]) begin
          $fwrite(f, "Register (27,6) Value: %h\n", PRED27_6_buffer[clk]);
        end
        if (PRED27_7_buffer[clk] != PRED27_7_buffer[!clk]) begin
          $fwrite(f, "Register (27,7) Value: %h\n", PRED27_7_buffer[clk]);
        end
        if (PRED27_8_buffer[clk] != PRED27_8_buffer[!clk]) begin
          $fwrite(f, "Register (27,8) Value: %h\n", PRED27_8_buffer[clk]);
        end
        if (PRED27_9_buffer[clk] != PRED27_9_buffer[!clk]) begin
          $fwrite(f, "Register (27,9) Value: %h\n", PRED27_9_buffer[clk]);
        end
        if (PRED27_10_buffer[clk] != PRED27_10_buffer[!clk]) begin
          $fwrite(f, "Register (27,10) Value: %h\n", PRED27_10_buffer[clk]);
        end
        if (PRED27_11_buffer[clk] != PRED27_11_buffer[!clk]) begin
          $fwrite(f, "Register (27,11) Value: %h\n", PRED27_11_buffer[clk]);
        end
        if (PRED27_12_buffer[clk] != PRED27_12_buffer[!clk]) begin
          $fwrite(f, "Register (27,12) Value: %h\n", PRED27_12_buffer[clk]);
        end
        if (PRED27_13_buffer[clk] != PRED27_13_buffer[!clk]) begin
          $fwrite(f, "Register (27,13) Value: %h\n", PRED27_13_buffer[clk]);
        end
        if (PRED27_14_buffer[clk] != PRED27_14_buffer[!clk]) begin
          $fwrite(f, "Register (27,14) Value: %h\n", PRED27_14_buffer[clk]);
        end
        if (PRED27_15_buffer[clk] != PRED27_15_buffer[!clk]) begin
          $fwrite(f, "Register (27,15) Value: %h\n", PRED27_15_buffer[clk]);
        end
        if (PRED27_16_buffer[clk] != PRED27_16_buffer[!clk]) begin
          $fwrite(f, "Register (27,16) Value: %h\n", PRED27_16_buffer[clk]);
        end
        if (PRED27_17_buffer[clk] != PRED27_17_buffer[!clk]) begin
          $fwrite(f, "Register (27,17) Value: %h\n", PRED27_17_buffer[clk]);
        end
        if (PRED27_18_buffer[clk] != PRED27_18_buffer[!clk]) begin
          $fwrite(f, "Register (27,18) Value: %h\n", PRED27_18_buffer[clk]);
        end
        if (PRED27_19_buffer[clk] != PRED27_19_buffer[!clk]) begin
          $fwrite(f, "Register (27,19) Value: %h\n", PRED27_19_buffer[clk]);
        end
        if (PRED27_20_buffer[clk] != PRED27_20_buffer[!clk]) begin
          $fwrite(f, "Register (27,20) Value: %h\n", PRED27_20_buffer[clk]);
        end
        if (PRED27_21_buffer[clk] != PRED27_21_buffer[!clk]) begin
          $fwrite(f, "Register (27,21) Value: %h\n", PRED27_21_buffer[clk]);
        end
        if (PRED27_22_buffer[clk] != PRED27_22_buffer[!clk]) begin
          $fwrite(f, "Register (27,22) Value: %h\n", PRED27_22_buffer[clk]);
        end
        if (PRED27_23_buffer[clk] != PRED27_23_buffer[!clk]) begin
          $fwrite(f, "Register (27,23) Value: %h\n", PRED27_23_buffer[clk]);
        end
        if (PRED27_24_buffer[clk] != PRED27_24_buffer[!clk]) begin
          $fwrite(f, "Register (27,24) Value: %h\n", PRED27_24_buffer[clk]);
        end
        if (PRED27_25_buffer[clk] != PRED27_25_buffer[!clk]) begin
          $fwrite(f, "Register (27,25) Value: %h\n", PRED27_25_buffer[clk]);
        end
        if (PRED27_26_buffer[clk] != PRED27_26_buffer[!clk]) begin
          $fwrite(f, "Register (27,26) Value: %h\n", PRED27_26_buffer[clk]);
        end
        if (PRED27_27_buffer[clk] != PRED27_27_buffer[!clk]) begin
          $fwrite(f, "Register (27,27) Value: %h\n", PRED27_27_buffer[clk]);
        end
        if (PRED27_28_buffer[clk] != PRED27_28_buffer[!clk]) begin
          $fwrite(f, "Register (27,28) Value: %h\n", PRED27_28_buffer[clk]);
        end
        if (PRED27_29_buffer[clk] != PRED27_29_buffer[!clk]) begin
          $fwrite(f, "Register (27,29) Value: %h\n", PRED27_29_buffer[clk]);
        end
        if (PRED27_30_buffer[clk] != PRED27_30_buffer[!clk]) begin
          $fwrite(f, "Register (27,30) Value: %h\n", PRED27_30_buffer[clk]);
        end
        if (PRED27_31_buffer[clk] != PRED27_31_buffer[!clk]) begin
          $fwrite(f, "Register (27,31) Value: %h\n", PRED27_31_buffer[clk]);
        end
        if (PRED28_0_buffer[clk] != PRED28_0_buffer[!clk]) begin
          $fwrite(f, "Register (28,0) Value: %h\n", PRED28_0_buffer[clk]);
        end
        if (PRED28_1_buffer[clk] != PRED28_1_buffer[!clk]) begin
          $fwrite(f, "Register (28,1) Value: %h\n", PRED28_1_buffer[clk]);
        end
        if (PRED28_2_buffer[clk] != PRED28_2_buffer[!clk]) begin
          $fwrite(f, "Register (28,2) Value: %h\n", PRED28_2_buffer[clk]);
        end
        if (PRED28_3_buffer[clk] != PRED28_3_buffer[!clk]) begin
          $fwrite(f, "Register (28,3) Value: %h\n", PRED28_3_buffer[clk]);
        end
        if (PRED28_4_buffer[clk] != PRED28_4_buffer[!clk]) begin
          $fwrite(f, "Register (28,4) Value: %h\n", PRED28_4_buffer[clk]);
        end
        if (PRED28_5_buffer[clk] != PRED28_5_buffer[!clk]) begin
          $fwrite(f, "Register (28,5) Value: %h\n", PRED28_5_buffer[clk]);
        end
        if (PRED28_6_buffer[clk] != PRED28_6_buffer[!clk]) begin
          $fwrite(f, "Register (28,6) Value: %h\n", PRED28_6_buffer[clk]);
        end
        if (PRED28_7_buffer[clk] != PRED28_7_buffer[!clk]) begin
          $fwrite(f, "Register (28,7) Value: %h\n", PRED28_7_buffer[clk]);
        end
        if (PRED28_8_buffer[clk] != PRED28_8_buffer[!clk]) begin
          $fwrite(f, "Register (28,8) Value: %h\n", PRED28_8_buffer[clk]);
        end
        if (PRED28_9_buffer[clk] != PRED28_9_buffer[!clk]) begin
          $fwrite(f, "Register (28,9) Value: %h\n", PRED28_9_buffer[clk]);
        end
        if (PRED28_10_buffer[clk] != PRED28_10_buffer[!clk]) begin
          $fwrite(f, "Register (28,10) Value: %h\n", PRED28_10_buffer[clk]);
        end
        if (PRED28_11_buffer[clk] != PRED28_11_buffer[!clk]) begin
          $fwrite(f, "Register (28,11) Value: %h\n", PRED28_11_buffer[clk]);
        end
        if (PRED28_12_buffer[clk] != PRED28_12_buffer[!clk]) begin
          $fwrite(f, "Register (28,12) Value: %h\n", PRED28_12_buffer[clk]);
        end
        if (PRED28_13_buffer[clk] != PRED28_13_buffer[!clk]) begin
          $fwrite(f, "Register (28,13) Value: %h\n", PRED28_13_buffer[clk]);
        end
        if (PRED28_14_buffer[clk] != PRED28_14_buffer[!clk]) begin
          $fwrite(f, "Register (28,14) Value: %h\n", PRED28_14_buffer[clk]);
        end
        if (PRED28_15_buffer[clk] != PRED28_15_buffer[!clk]) begin
          $fwrite(f, "Register (28,15) Value: %h\n", PRED28_15_buffer[clk]);
        end
        if (PRED28_16_buffer[clk] != PRED28_16_buffer[!clk]) begin
          $fwrite(f, "Register (28,16) Value: %h\n", PRED28_16_buffer[clk]);
        end
        if (PRED28_17_buffer[clk] != PRED28_17_buffer[!clk]) begin
          $fwrite(f, "Register (28,17) Value: %h\n", PRED28_17_buffer[clk]);
        end
        if (PRED28_18_buffer[clk] != PRED28_18_buffer[!clk]) begin
          $fwrite(f, "Register (28,18) Value: %h\n", PRED28_18_buffer[clk]);
        end
        if (PRED28_19_buffer[clk] != PRED28_19_buffer[!clk]) begin
          $fwrite(f, "Register (28,19) Value: %h\n", PRED28_19_buffer[clk]);
        end
        if (PRED28_20_buffer[clk] != PRED28_20_buffer[!clk]) begin
          $fwrite(f, "Register (28,20) Value: %h\n", PRED28_20_buffer[clk]);
        end
        if (PRED28_21_buffer[clk] != PRED28_21_buffer[!clk]) begin
          $fwrite(f, "Register (28,21) Value: %h\n", PRED28_21_buffer[clk]);
        end
        if (PRED28_22_buffer[clk] != PRED28_22_buffer[!clk]) begin
          $fwrite(f, "Register (28,22) Value: %h\n", PRED28_22_buffer[clk]);
        end
        if (PRED28_23_buffer[clk] != PRED28_23_buffer[!clk]) begin
          $fwrite(f, "Register (28,23) Value: %h\n", PRED28_23_buffer[clk]);
        end
        if (PRED28_24_buffer[clk] != PRED28_24_buffer[!clk]) begin
          $fwrite(f, "Register (28,24) Value: %h\n", PRED28_24_buffer[clk]);
        end
        if (PRED28_25_buffer[clk] != PRED28_25_buffer[!clk]) begin
          $fwrite(f, "Register (28,25) Value: %h\n", PRED28_25_buffer[clk]);
        end
        if (PRED28_26_buffer[clk] != PRED28_26_buffer[!clk]) begin
          $fwrite(f, "Register (28,26) Value: %h\n", PRED28_26_buffer[clk]);
        end
        if (PRED28_27_buffer[clk] != PRED28_27_buffer[!clk]) begin
          $fwrite(f, "Register (28,27) Value: %h\n", PRED28_27_buffer[clk]);
        end
        if (PRED28_28_buffer[clk] != PRED28_28_buffer[!clk]) begin
          $fwrite(f, "Register (28,28) Value: %h\n", PRED28_28_buffer[clk]);
        end
        if (PRED28_29_buffer[clk] != PRED28_29_buffer[!clk]) begin
          $fwrite(f, "Register (28,29) Value: %h\n", PRED28_29_buffer[clk]);
        end
        if (PRED28_30_buffer[clk] != PRED28_30_buffer[!clk]) begin
          $fwrite(f, "Register (28,30) Value: %h\n", PRED28_30_buffer[clk]);
        end
        if (PRED28_31_buffer[clk] != PRED28_31_buffer[!clk]) begin
          $fwrite(f, "Register (28,31) Value: %h\n", PRED28_31_buffer[clk]);
        end
        if (PRED29_0_buffer[clk] != PRED29_0_buffer[!clk]) begin
          $fwrite(f, "Register (29,0) Value: %h\n", PRED29_0_buffer[clk]);
        end
        if (PRED29_1_buffer[clk] != PRED29_1_buffer[!clk]) begin
          $fwrite(f, "Register (29,1) Value: %h\n", PRED29_1_buffer[clk]);
        end
        if (PRED29_2_buffer[clk] != PRED29_2_buffer[!clk]) begin
          $fwrite(f, "Register (29,2) Value: %h\n", PRED29_2_buffer[clk]);
        end
        if (PRED29_3_buffer[clk] != PRED29_3_buffer[!clk]) begin
          $fwrite(f, "Register (29,3) Value: %h\n", PRED29_3_buffer[clk]);
        end
        if (PRED29_4_buffer[clk] != PRED29_4_buffer[!clk]) begin
          $fwrite(f, "Register (29,4) Value: %h\n", PRED29_4_buffer[clk]);
        end
        if (PRED29_5_buffer[clk] != PRED29_5_buffer[!clk]) begin
          $fwrite(f, "Register (29,5) Value: %h\n", PRED29_5_buffer[clk]);
        end
        if (PRED29_6_buffer[clk] != PRED29_6_buffer[!clk]) begin
          $fwrite(f, "Register (29,6) Value: %h\n", PRED29_6_buffer[clk]);
        end
        if (PRED29_7_buffer[clk] != PRED29_7_buffer[!clk]) begin
          $fwrite(f, "Register (29,7) Value: %h\n", PRED29_7_buffer[clk]);
        end
        if (PRED29_8_buffer[clk] != PRED29_8_buffer[!clk]) begin
          $fwrite(f, "Register (29,8) Value: %h\n", PRED29_8_buffer[clk]);
        end
        if (PRED29_9_buffer[clk] != PRED29_9_buffer[!clk]) begin
          $fwrite(f, "Register (29,9) Value: %h\n", PRED29_9_buffer[clk]);
        end
        if (PRED29_10_buffer[clk] != PRED29_10_buffer[!clk]) begin
          $fwrite(f, "Register (29,10) Value: %h\n", PRED29_10_buffer[clk]);
        end
        if (PRED29_11_buffer[clk] != PRED29_11_buffer[!clk]) begin
          $fwrite(f, "Register (29,11) Value: %h\n", PRED29_11_buffer[clk]);
        end
        if (PRED29_12_buffer[clk] != PRED29_12_buffer[!clk]) begin
          $fwrite(f, "Register (29,12) Value: %h\n", PRED29_12_buffer[clk]);
        end
        if (PRED29_13_buffer[clk] != PRED29_13_buffer[!clk]) begin
          $fwrite(f, "Register (29,13) Value: %h\n", PRED29_13_buffer[clk]);
        end
        if (PRED29_14_buffer[clk] != PRED29_14_buffer[!clk]) begin
          $fwrite(f, "Register (29,14) Value: %h\n", PRED29_14_buffer[clk]);
        end
        if (PRED29_15_buffer[clk] != PRED29_15_buffer[!clk]) begin
          $fwrite(f, "Register (29,15) Value: %h\n", PRED29_15_buffer[clk]);
        end
        if (PRED29_16_buffer[clk] != PRED29_16_buffer[!clk]) begin
          $fwrite(f, "Register (29,16) Value: %h\n", PRED29_16_buffer[clk]);
        end
        if (PRED29_17_buffer[clk] != PRED29_17_buffer[!clk]) begin
          $fwrite(f, "Register (29,17) Value: %h\n", PRED29_17_buffer[clk]);
        end
        if (PRED29_18_buffer[clk] != PRED29_18_buffer[!clk]) begin
          $fwrite(f, "Register (29,18) Value: %h\n", PRED29_18_buffer[clk]);
        end
        if (PRED29_19_buffer[clk] != PRED29_19_buffer[!clk]) begin
          $fwrite(f, "Register (29,19) Value: %h\n", PRED29_19_buffer[clk]);
        end
        if (PRED29_20_buffer[clk] != PRED29_20_buffer[!clk]) begin
          $fwrite(f, "Register (29,20) Value: %h\n", PRED29_20_buffer[clk]);
        end
        if (PRED29_21_buffer[clk] != PRED29_21_buffer[!clk]) begin
          $fwrite(f, "Register (29,21) Value: %h\n", PRED29_21_buffer[clk]);
        end
        if (PRED29_22_buffer[clk] != PRED29_22_buffer[!clk]) begin
          $fwrite(f, "Register (29,22) Value: %h\n", PRED29_22_buffer[clk]);
        end
        if (PRED29_23_buffer[clk] != PRED29_23_buffer[!clk]) begin
          $fwrite(f, "Register (29,23) Value: %h\n", PRED29_23_buffer[clk]);
        end
        if (PRED29_24_buffer[clk] != PRED29_24_buffer[!clk]) begin
          $fwrite(f, "Register (29,24) Value: %h\n", PRED29_24_buffer[clk]);
        end
        if (PRED29_25_buffer[clk] != PRED29_25_buffer[!clk]) begin
          $fwrite(f, "Register (29,25) Value: %h\n", PRED29_25_buffer[clk]);
        end
        if (PRED29_26_buffer[clk] != PRED29_26_buffer[!clk]) begin
          $fwrite(f, "Register (29,26) Value: %h\n", PRED29_26_buffer[clk]);
        end
        if (PRED29_27_buffer[clk] != PRED29_27_buffer[!clk]) begin
          $fwrite(f, "Register (29,27) Value: %h\n", PRED29_27_buffer[clk]);
        end
        if (PRED29_28_buffer[clk] != PRED29_28_buffer[!clk]) begin
          $fwrite(f, "Register (29,28) Value: %h\n", PRED29_28_buffer[clk]);
        end
        if (PRED29_29_buffer[clk] != PRED29_29_buffer[!clk]) begin
          $fwrite(f, "Register (29,29) Value: %h\n", PRED29_29_buffer[clk]);
        end
        if (PRED29_30_buffer[clk] != PRED29_30_buffer[!clk]) begin
          $fwrite(f, "Register (29,30) Value: %h\n", PRED29_30_buffer[clk]);
        end
        if (PRED29_31_buffer[clk] != PRED29_31_buffer[!clk]) begin
          $fwrite(f, "Register (29,31) Value: %h\n", PRED29_31_buffer[clk]);
        end
        if (PRED30_0_buffer[clk] != PRED30_0_buffer[!clk]) begin
          $fwrite(f, "Register (30,0) Value: %h\n", PRED30_0_buffer[clk]);
        end
        if (PRED30_1_buffer[clk] != PRED30_1_buffer[!clk]) begin
          $fwrite(f, "Register (30,1) Value: %h\n", PRED30_1_buffer[clk]);
        end
        if (PRED30_2_buffer[clk] != PRED30_2_buffer[!clk]) begin
          $fwrite(f, "Register (30,2) Value: %h\n", PRED30_2_buffer[clk]);
        end
        if (PRED30_3_buffer[clk] != PRED30_3_buffer[!clk]) begin
          $fwrite(f, "Register (30,3) Value: %h\n", PRED30_3_buffer[clk]);
        end
        if (PRED30_4_buffer[clk] != PRED30_4_buffer[!clk]) begin
          $fwrite(f, "Register (30,4) Value: %h\n", PRED30_4_buffer[clk]);
        end
        if (PRED30_5_buffer[clk] != PRED30_5_buffer[!clk]) begin
          $fwrite(f, "Register (30,5) Value: %h\n", PRED30_5_buffer[clk]);
        end
        if (PRED30_6_buffer[clk] != PRED30_6_buffer[!clk]) begin
          $fwrite(f, "Register (30,6) Value: %h\n", PRED30_6_buffer[clk]);
        end
        if (PRED30_7_buffer[clk] != PRED30_7_buffer[!clk]) begin
          $fwrite(f, "Register (30,7) Value: %h\n", PRED30_7_buffer[clk]);
        end
        if (PRED30_8_buffer[clk] != PRED30_8_buffer[!clk]) begin
          $fwrite(f, "Register (30,8) Value: %h\n", PRED30_8_buffer[clk]);
        end
        if (PRED30_9_buffer[clk] != PRED30_9_buffer[!clk]) begin
          $fwrite(f, "Register (30,9) Value: %h\n", PRED30_9_buffer[clk]);
        end
        if (PRED30_10_buffer[clk] != PRED30_10_buffer[!clk]) begin
          $fwrite(f, "Register (30,10) Value: %h\n", PRED30_10_buffer[clk]);
        end
        if (PRED30_11_buffer[clk] != PRED30_11_buffer[!clk]) begin
          $fwrite(f, "Register (30,11) Value: %h\n", PRED30_11_buffer[clk]);
        end
        if (PRED30_12_buffer[clk] != PRED30_12_buffer[!clk]) begin
          $fwrite(f, "Register (30,12) Value: %h\n", PRED30_12_buffer[clk]);
        end
        if (PRED30_13_buffer[clk] != PRED30_13_buffer[!clk]) begin
          $fwrite(f, "Register (30,13) Value: %h\n", PRED30_13_buffer[clk]);
        end
        if (PRED30_14_buffer[clk] != PRED30_14_buffer[!clk]) begin
          $fwrite(f, "Register (30,14) Value: %h\n", PRED30_14_buffer[clk]);
        end
        if (PRED30_15_buffer[clk] != PRED30_15_buffer[!clk]) begin
          $fwrite(f, "Register (30,15) Value: %h\n", PRED30_15_buffer[clk]);
        end
        if (PRED30_16_buffer[clk] != PRED30_16_buffer[!clk]) begin
          $fwrite(f, "Register (30,16) Value: %h\n", PRED30_16_buffer[clk]);
        end
        if (PRED30_17_buffer[clk] != PRED30_17_buffer[!clk]) begin
          $fwrite(f, "Register (30,17) Value: %h\n", PRED30_17_buffer[clk]);
        end
        if (PRED30_18_buffer[clk] != PRED30_18_buffer[!clk]) begin
          $fwrite(f, "Register (30,18) Value: %h\n", PRED30_18_buffer[clk]);
        end
        if (PRED30_19_buffer[clk] != PRED30_19_buffer[!clk]) begin
          $fwrite(f, "Register (30,19) Value: %h\n", PRED30_19_buffer[clk]);
        end
        if (PRED30_20_buffer[clk] != PRED30_20_buffer[!clk]) begin
          $fwrite(f, "Register (30,20) Value: %h\n", PRED30_20_buffer[clk]);
        end
        if (PRED30_21_buffer[clk] != PRED30_21_buffer[!clk]) begin
          $fwrite(f, "Register (30,21) Value: %h\n", PRED30_21_buffer[clk]);
        end
        if (PRED30_22_buffer[clk] != PRED30_22_buffer[!clk]) begin
          $fwrite(f, "Register (30,22) Value: %h\n", PRED30_22_buffer[clk]);
        end
        if (PRED30_23_buffer[clk] != PRED30_23_buffer[!clk]) begin
          $fwrite(f, "Register (30,23) Value: %h\n", PRED30_23_buffer[clk]);
        end
        if (PRED30_24_buffer[clk] != PRED30_24_buffer[!clk]) begin
          $fwrite(f, "Register (30,24) Value: %h\n", PRED30_24_buffer[clk]);
        end
        if (PRED30_25_buffer[clk] != PRED30_25_buffer[!clk]) begin
          $fwrite(f, "Register (30,25) Value: %h\n", PRED30_25_buffer[clk]);
        end
        if (PRED30_26_buffer[clk] != PRED30_26_buffer[!clk]) begin
          $fwrite(f, "Register (30,26) Value: %h\n", PRED30_26_buffer[clk]);
        end
        if (PRED30_27_buffer[clk] != PRED30_27_buffer[!clk]) begin
          $fwrite(f, "Register (30,27) Value: %h\n", PRED30_27_buffer[clk]);
        end
        if (PRED30_28_buffer[clk] != PRED30_28_buffer[!clk]) begin
          $fwrite(f, "Register (30,28) Value: %h\n", PRED30_28_buffer[clk]);
        end
        if (PRED30_29_buffer[clk] != PRED30_29_buffer[!clk]) begin
          $fwrite(f, "Register (30,29) Value: %h\n", PRED30_29_buffer[clk]);
        end
        if (PRED30_30_buffer[clk] != PRED30_30_buffer[!clk]) begin
          $fwrite(f, "Register (30,30) Value: %h\n", PRED30_30_buffer[clk]);
        end
        if (PRED30_31_buffer[clk] != PRED30_31_buffer[!clk]) begin
          $fwrite(f, "Register (30,31) Value: %h\n", PRED30_31_buffer[clk]);
        end
        if (PRED31_0_buffer[clk] != PRED31_0_buffer[!clk]) begin
          $fwrite(f, "Register (31,0) Value: %h\n", PRED31_0_buffer[clk]);
        end
        if (PRED31_1_buffer[clk] != PRED31_1_buffer[!clk]) begin
          $fwrite(f, "Register (31,1) Value: %h\n", PRED31_1_buffer[clk]);
        end
        if (PRED31_2_buffer[clk] != PRED31_2_buffer[!clk]) begin
          $fwrite(f, "Register (31,2) Value: %h\n", PRED31_2_buffer[clk]);
        end
        if (PRED31_3_buffer[clk] != PRED31_3_buffer[!clk]) begin
          $fwrite(f, "Register (31,3) Value: %h\n", PRED31_3_buffer[clk]);
        end
        if (PRED31_4_buffer[clk] != PRED31_4_buffer[!clk]) begin
          $fwrite(f, "Register (31,4) Value: %h\n", PRED31_4_buffer[clk]);
        end
        if (PRED31_5_buffer[clk] != PRED31_5_buffer[!clk]) begin
          $fwrite(f, "Register (31,5) Value: %h\n", PRED31_5_buffer[clk]);
        end
        if (PRED31_6_buffer[clk] != PRED31_6_buffer[!clk]) begin
          $fwrite(f, "Register (31,6) Value: %h\n", PRED31_6_buffer[clk]);
        end
        if (PRED31_7_buffer[clk] != PRED31_7_buffer[!clk]) begin
          $fwrite(f, "Register (31,7) Value: %h\n", PRED31_7_buffer[clk]);
        end
        if (PRED31_8_buffer[clk] != PRED31_8_buffer[!clk]) begin
          $fwrite(f, "Register (31,8) Value: %h\n", PRED31_8_buffer[clk]);
        end
        if (PRED31_9_buffer[clk] != PRED31_9_buffer[!clk]) begin
          $fwrite(f, "Register (31,9) Value: %h\n", PRED31_9_buffer[clk]);
        end
        if (PRED31_10_buffer[clk] != PRED31_10_buffer[!clk]) begin
          $fwrite(f, "Register (31,10) Value: %h\n", PRED31_10_buffer[clk]);
        end
        if (PRED31_11_buffer[clk] != PRED31_11_buffer[!clk]) begin
          $fwrite(f, "Register (31,11) Value: %h\n", PRED31_11_buffer[clk]);
        end
        if (PRED31_12_buffer[clk] != PRED31_12_buffer[!clk]) begin
          $fwrite(f, "Register (31,12) Value: %h\n", PRED31_12_buffer[clk]);
        end
        if (PRED31_13_buffer[clk] != PRED31_13_buffer[!clk]) begin
          $fwrite(f, "Register (31,13) Value: %h\n", PRED31_13_buffer[clk]);
        end
        if (PRED31_14_buffer[clk] != PRED31_14_buffer[!clk]) begin
          $fwrite(f, "Register (31,14) Value: %h\n", PRED31_14_buffer[clk]);
        end
        if (PRED31_15_buffer[clk] != PRED31_15_buffer[!clk]) begin
          $fwrite(f, "Register (31,15) Value: %h\n", PRED31_15_buffer[clk]);
        end
        if (PRED31_16_buffer[clk] != PRED31_16_buffer[!clk]) begin
          $fwrite(f, "Register (31,16) Value: %h\n", PRED31_16_buffer[clk]);
        end
        if (PRED31_17_buffer[clk] != PRED31_17_buffer[!clk]) begin
          $fwrite(f, "Register (31,17) Value: %h\n", PRED31_17_buffer[clk]);
        end
        if (PRED31_18_buffer[clk] != PRED31_18_buffer[!clk]) begin
          $fwrite(f, "Register (31,18) Value: %h\n", PRED31_18_buffer[clk]);
        end
        if (PRED31_19_buffer[clk] != PRED31_19_buffer[!clk]) begin
          $fwrite(f, "Register (31,19) Value: %h\n", PRED31_19_buffer[clk]);
        end
        if (PRED31_20_buffer[clk] != PRED31_20_buffer[!clk]) begin
          $fwrite(f, "Register (31,20) Value: %h\n", PRED31_20_buffer[clk]);
        end
        if (PRED31_21_buffer[clk] != PRED31_21_buffer[!clk]) begin
          $fwrite(f, "Register (31,21) Value: %h\n", PRED31_21_buffer[clk]);
        end
        if (PRED31_22_buffer[clk] != PRED31_22_buffer[!clk]) begin
          $fwrite(f, "Register (31,22) Value: %h\n", PRED31_22_buffer[clk]);
        end
        if (PRED31_23_buffer[clk] != PRED31_23_buffer[!clk]) begin
          $fwrite(f, "Register (31,23) Value: %h\n", PRED31_23_buffer[clk]);
        end
        if (PRED31_24_buffer[clk] != PRED31_24_buffer[!clk]) begin
          $fwrite(f, "Register (31,24) Value: %h\n", PRED31_24_buffer[clk]);
        end
        if (PRED31_25_buffer[clk] != PRED31_25_buffer[!clk]) begin
          $fwrite(f, "Register (31,25) Value: %h\n", PRED31_25_buffer[clk]);
        end
        if (PRED31_26_buffer[clk] != PRED31_26_buffer[!clk]) begin
          $fwrite(f, "Register (31,26) Value: %h\n", PRED31_26_buffer[clk]);
        end
        if (PRED31_27_buffer[clk] != PRED31_27_buffer[!clk]) begin
          $fwrite(f, "Register (31,27) Value: %h\n", PRED31_27_buffer[clk]);
        end
        if (PRED31_28_buffer[clk] != PRED31_28_buffer[!clk]) begin
          $fwrite(f, "Register (31,28) Value: %h\n", PRED31_28_buffer[clk]);
        end
        if (PRED31_29_buffer[clk] != PRED31_29_buffer[!clk]) begin
          $fwrite(f, "Register (31,29) Value: %h\n", PRED31_29_buffer[clk]);
        end
        if (PRED31_30_buffer[clk] != PRED31_30_buffer[!clk]) begin
          $fwrite(f, "Register (31,30) Value: %h\n", PRED31_30_buffer[clk]);
        end
        if (PRED31_31_buffer[clk] != PRED31_31_buffer[!clk]) begin
          $fwrite(f, "Register (31,31) Value: %h\n", PRED31_31_buffer[clk]);
        end
        if (PRED32_0_buffer[clk] != PRED32_0_buffer[!clk]) begin
          $fwrite(f, "Register (32,0) Value: %h\n", PRED32_0_buffer[clk]);
        end
        if (PRED32_1_buffer[clk] != PRED32_1_buffer[!clk]) begin
          $fwrite(f, "Register (32,1) Value: %h\n", PRED32_1_buffer[clk]);
        end
        if (PRED32_2_buffer[clk] != PRED32_2_buffer[!clk]) begin
          $fwrite(f, "Register (32,2) Value: %h\n", PRED32_2_buffer[clk]);
        end
        if (PRED32_3_buffer[clk] != PRED32_3_buffer[!clk]) begin
          $fwrite(f, "Register (32,3) Value: %h\n", PRED32_3_buffer[clk]);
        end
        if (PRED32_4_buffer[clk] != PRED32_4_buffer[!clk]) begin
          $fwrite(f, "Register (32,4) Value: %h\n", PRED32_4_buffer[clk]);
        end
        if (PRED32_5_buffer[clk] != PRED32_5_buffer[!clk]) begin
          $fwrite(f, "Register (32,5) Value: %h\n", PRED32_5_buffer[clk]);
        end
        if (PRED32_6_buffer[clk] != PRED32_6_buffer[!clk]) begin
          $fwrite(f, "Register (32,6) Value: %h\n", PRED32_6_buffer[clk]);
        end
        if (PRED32_7_buffer[clk] != PRED32_7_buffer[!clk]) begin
          $fwrite(f, "Register (32,7) Value: %h\n", PRED32_7_buffer[clk]);
        end
        if (PRED32_8_buffer[clk] != PRED32_8_buffer[!clk]) begin
          $fwrite(f, "Register (32,8) Value: %h\n", PRED32_8_buffer[clk]);
        end
        if (PRED32_9_buffer[clk] != PRED32_9_buffer[!clk]) begin
          $fwrite(f, "Register (32,9) Value: %h\n", PRED32_9_buffer[clk]);
        end
        if (PRED32_10_buffer[clk] != PRED32_10_buffer[!clk]) begin
          $fwrite(f, "Register (32,10) Value: %h\n", PRED32_10_buffer[clk]);
        end
        if (PRED32_11_buffer[clk] != PRED32_11_buffer[!clk]) begin
          $fwrite(f, "Register (32,11) Value: %h\n", PRED32_11_buffer[clk]);
        end
        if (PRED32_12_buffer[clk] != PRED32_12_buffer[!clk]) begin
          $fwrite(f, "Register (32,12) Value: %h\n", PRED32_12_buffer[clk]);
        end
        if (PRED32_13_buffer[clk] != PRED32_13_buffer[!clk]) begin
          $fwrite(f, "Register (32,13) Value: %h\n", PRED32_13_buffer[clk]);
        end
        if (PRED32_14_buffer[clk] != PRED32_14_buffer[!clk]) begin
          $fwrite(f, "Register (32,14) Value: %h\n", PRED32_14_buffer[clk]);
        end
        if (PRED32_15_buffer[clk] != PRED32_15_buffer[!clk]) begin
          $fwrite(f, "Register (32,15) Value: %h\n", PRED32_15_buffer[clk]);
        end
        if (PRED32_16_buffer[clk] != PRED32_16_buffer[!clk]) begin
          $fwrite(f, "Register (32,16) Value: %h\n", PRED32_16_buffer[clk]);
        end
        if (PRED32_17_buffer[clk] != PRED32_17_buffer[!clk]) begin
          $fwrite(f, "Register (32,17) Value: %h\n", PRED32_17_buffer[clk]);
        end
        if (PRED32_18_buffer[clk] != PRED32_18_buffer[!clk]) begin
          $fwrite(f, "Register (32,18) Value: %h\n", PRED32_18_buffer[clk]);
        end
        if (PRED32_19_buffer[clk] != PRED32_19_buffer[!clk]) begin
          $fwrite(f, "Register (32,19) Value: %h\n", PRED32_19_buffer[clk]);
        end
        if (PRED32_20_buffer[clk] != PRED32_20_buffer[!clk]) begin
          $fwrite(f, "Register (32,20) Value: %h\n", PRED32_20_buffer[clk]);
        end
        if (PRED32_21_buffer[clk] != PRED32_21_buffer[!clk]) begin
          $fwrite(f, "Register (32,21) Value: %h\n", PRED32_21_buffer[clk]);
        end
        if (PRED32_22_buffer[clk] != PRED32_22_buffer[!clk]) begin
          $fwrite(f, "Register (32,22) Value: %h\n", PRED32_22_buffer[clk]);
        end
        if (PRED32_23_buffer[clk] != PRED32_23_buffer[!clk]) begin
          $fwrite(f, "Register (32,23) Value: %h\n", PRED32_23_buffer[clk]);
        end
        if (PRED32_24_buffer[clk] != PRED32_24_buffer[!clk]) begin
          $fwrite(f, "Register (32,24) Value: %h\n", PRED32_24_buffer[clk]);
        end
        if (PRED32_25_buffer[clk] != PRED32_25_buffer[!clk]) begin
          $fwrite(f, "Register (32,25) Value: %h\n", PRED32_25_buffer[clk]);
        end
        if (PRED32_26_buffer[clk] != PRED32_26_buffer[!clk]) begin
          $fwrite(f, "Register (32,26) Value: %h\n", PRED32_26_buffer[clk]);
        end
        if (PRED32_27_buffer[clk] != PRED32_27_buffer[!clk]) begin
          $fwrite(f, "Register (32,27) Value: %h\n", PRED32_27_buffer[clk]);
        end
        if (PRED32_28_buffer[clk] != PRED32_28_buffer[!clk]) begin
          $fwrite(f, "Register (32,28) Value: %h\n", PRED32_28_buffer[clk]);
        end
        if (PRED32_29_buffer[clk] != PRED32_29_buffer[!clk]) begin
          $fwrite(f, "Register (32,29) Value: %h\n", PRED32_29_buffer[clk]);
        end
        if (PRED32_30_buffer[clk] != PRED32_30_buffer[!clk]) begin
          $fwrite(f, "Register (32,30) Value: %h\n", PRED32_30_buffer[clk]);
        end
        if (PRED32_31_buffer[clk] != PRED32_31_buffer[!clk]) begin
          $fwrite(f, "Register (32,31) Value: %h\n", PRED32_31_buffer[clk]);
        end
        if (PRED33_0_buffer[clk] != PRED33_0_buffer[!clk]) begin
          $fwrite(f, "Register (33,0) Value: %h\n", PRED33_0_buffer[clk]);
        end
        if (PRED33_1_buffer[clk] != PRED33_1_buffer[!clk]) begin
          $fwrite(f, "Register (33,1) Value: %h\n", PRED33_1_buffer[clk]);
        end
        if (PRED33_2_buffer[clk] != PRED33_2_buffer[!clk]) begin
          $fwrite(f, "Register (33,2) Value: %h\n", PRED33_2_buffer[clk]);
        end
        if (PRED33_3_buffer[clk] != PRED33_3_buffer[!clk]) begin
          $fwrite(f, "Register (33,3) Value: %h\n", PRED33_3_buffer[clk]);
        end
        if (PRED33_4_buffer[clk] != PRED33_4_buffer[!clk]) begin
          $fwrite(f, "Register (33,4) Value: %h\n", PRED33_4_buffer[clk]);
        end
        if (PRED33_5_buffer[clk] != PRED33_5_buffer[!clk]) begin
          $fwrite(f, "Register (33,5) Value: %h\n", PRED33_5_buffer[clk]);
        end
        if (PRED33_6_buffer[clk] != PRED33_6_buffer[!clk]) begin
          $fwrite(f, "Register (33,6) Value: %h\n", PRED33_6_buffer[clk]);
        end
        if (PRED33_7_buffer[clk] != PRED33_7_buffer[!clk]) begin
          $fwrite(f, "Register (33,7) Value: %h\n", PRED33_7_buffer[clk]);
        end
        if (PRED33_8_buffer[clk] != PRED33_8_buffer[!clk]) begin
          $fwrite(f, "Register (33,8) Value: %h\n", PRED33_8_buffer[clk]);
        end
        if (PRED33_9_buffer[clk] != PRED33_9_buffer[!clk]) begin
          $fwrite(f, "Register (33,9) Value: %h\n", PRED33_9_buffer[clk]);
        end
        if (PRED33_10_buffer[clk] != PRED33_10_buffer[!clk]) begin
          $fwrite(f, "Register (33,10) Value: %h\n", PRED33_10_buffer[clk]);
        end
        if (PRED33_11_buffer[clk] != PRED33_11_buffer[!clk]) begin
          $fwrite(f, "Register (33,11) Value: %h\n", PRED33_11_buffer[clk]);
        end
        if (PRED33_12_buffer[clk] != PRED33_12_buffer[!clk]) begin
          $fwrite(f, "Register (33,12) Value: %h\n", PRED33_12_buffer[clk]);
        end
        if (PRED33_13_buffer[clk] != PRED33_13_buffer[!clk]) begin
          $fwrite(f, "Register (33,13) Value: %h\n", PRED33_13_buffer[clk]);
        end
        if (PRED33_14_buffer[clk] != PRED33_14_buffer[!clk]) begin
          $fwrite(f, "Register (33,14) Value: %h\n", PRED33_14_buffer[clk]);
        end
        if (PRED33_15_buffer[clk] != PRED33_15_buffer[!clk]) begin
          $fwrite(f, "Register (33,15) Value: %h\n", PRED33_15_buffer[clk]);
        end
        if (PRED33_16_buffer[clk] != PRED33_16_buffer[!clk]) begin
          $fwrite(f, "Register (33,16) Value: %h\n", PRED33_16_buffer[clk]);
        end
        if (PRED33_17_buffer[clk] != PRED33_17_buffer[!clk]) begin
          $fwrite(f, "Register (33,17) Value: %h\n", PRED33_17_buffer[clk]);
        end
        if (PRED33_18_buffer[clk] != PRED33_18_buffer[!clk]) begin
          $fwrite(f, "Register (33,18) Value: %h\n", PRED33_18_buffer[clk]);
        end
        if (PRED33_19_buffer[clk] != PRED33_19_buffer[!clk]) begin
          $fwrite(f, "Register (33,19) Value: %h\n", PRED33_19_buffer[clk]);
        end
        if (PRED33_20_buffer[clk] != PRED33_20_buffer[!clk]) begin
          $fwrite(f, "Register (33,20) Value: %h\n", PRED33_20_buffer[clk]);
        end
        if (PRED33_21_buffer[clk] != PRED33_21_buffer[!clk]) begin
          $fwrite(f, "Register (33,21) Value: %h\n", PRED33_21_buffer[clk]);
        end
        if (PRED33_22_buffer[clk] != PRED33_22_buffer[!clk]) begin
          $fwrite(f, "Register (33,22) Value: %h\n", PRED33_22_buffer[clk]);
        end
        if (PRED33_23_buffer[clk] != PRED33_23_buffer[!clk]) begin
          $fwrite(f, "Register (33,23) Value: %h\n", PRED33_23_buffer[clk]);
        end
        if (PRED33_24_buffer[clk] != PRED33_24_buffer[!clk]) begin
          $fwrite(f, "Register (33,24) Value: %h\n", PRED33_24_buffer[clk]);
        end
        if (PRED33_25_buffer[clk] != PRED33_25_buffer[!clk]) begin
          $fwrite(f, "Register (33,25) Value: %h\n", PRED33_25_buffer[clk]);
        end
        if (PRED33_26_buffer[clk] != PRED33_26_buffer[!clk]) begin
          $fwrite(f, "Register (33,26) Value: %h\n", PRED33_26_buffer[clk]);
        end
        if (PRED33_27_buffer[clk] != PRED33_27_buffer[!clk]) begin
          $fwrite(f, "Register (33,27) Value: %h\n", PRED33_27_buffer[clk]);
        end
        if (PRED33_28_buffer[clk] != PRED33_28_buffer[!clk]) begin
          $fwrite(f, "Register (33,28) Value: %h\n", PRED33_28_buffer[clk]);
        end
        if (PRED33_29_buffer[clk] != PRED33_29_buffer[!clk]) begin
          $fwrite(f, "Register (33,29) Value: %h\n", PRED33_29_buffer[clk]);
        end
        if (PRED33_30_buffer[clk] != PRED33_30_buffer[!clk]) begin
          $fwrite(f, "Register (33,30) Value: %h\n", PRED33_30_buffer[clk]);
        end
        if (PRED33_31_buffer[clk] != PRED33_31_buffer[!clk]) begin
          $fwrite(f, "Register (33,31) Value: %h\n", PRED33_31_buffer[clk]);
        end
        if (PRED34_0_buffer[clk] != PRED34_0_buffer[!clk]) begin
          $fwrite(f, "Register (34,0) Value: %h\n", PRED34_0_buffer[clk]);
        end
        if (PRED34_1_buffer[clk] != PRED34_1_buffer[!clk]) begin
          $fwrite(f, "Register (34,1) Value: %h\n", PRED34_1_buffer[clk]);
        end
        if (PRED34_2_buffer[clk] != PRED34_2_buffer[!clk]) begin
          $fwrite(f, "Register (34,2) Value: %h\n", PRED34_2_buffer[clk]);
        end
        if (PRED34_3_buffer[clk] != PRED34_3_buffer[!clk]) begin
          $fwrite(f, "Register (34,3) Value: %h\n", PRED34_3_buffer[clk]);
        end
        if (PRED34_4_buffer[clk] != PRED34_4_buffer[!clk]) begin
          $fwrite(f, "Register (34,4) Value: %h\n", PRED34_4_buffer[clk]);
        end
        if (PRED34_5_buffer[clk] != PRED34_5_buffer[!clk]) begin
          $fwrite(f, "Register (34,5) Value: %h\n", PRED34_5_buffer[clk]);
        end
        if (PRED34_6_buffer[clk] != PRED34_6_buffer[!clk]) begin
          $fwrite(f, "Register (34,6) Value: %h\n", PRED34_6_buffer[clk]);
        end
        if (PRED34_7_buffer[clk] != PRED34_7_buffer[!clk]) begin
          $fwrite(f, "Register (34,7) Value: %h\n", PRED34_7_buffer[clk]);
        end
        if (PRED34_8_buffer[clk] != PRED34_8_buffer[!clk]) begin
          $fwrite(f, "Register (34,8) Value: %h\n", PRED34_8_buffer[clk]);
        end
        if (PRED34_9_buffer[clk] != PRED34_9_buffer[!clk]) begin
          $fwrite(f, "Register (34,9) Value: %h\n", PRED34_9_buffer[clk]);
        end
        if (PRED34_10_buffer[clk] != PRED34_10_buffer[!clk]) begin
          $fwrite(f, "Register (34,10) Value: %h\n", PRED34_10_buffer[clk]);
        end
        if (PRED34_11_buffer[clk] != PRED34_11_buffer[!clk]) begin
          $fwrite(f, "Register (34,11) Value: %h\n", PRED34_11_buffer[clk]);
        end
        if (PRED34_12_buffer[clk] != PRED34_12_buffer[!clk]) begin
          $fwrite(f, "Register (34,12) Value: %h\n", PRED34_12_buffer[clk]);
        end
        if (PRED34_13_buffer[clk] != PRED34_13_buffer[!clk]) begin
          $fwrite(f, "Register (34,13) Value: %h\n", PRED34_13_buffer[clk]);
        end
        if (PRED34_14_buffer[clk] != PRED34_14_buffer[!clk]) begin
          $fwrite(f, "Register (34,14) Value: %h\n", PRED34_14_buffer[clk]);
        end
        if (PRED34_15_buffer[clk] != PRED34_15_buffer[!clk]) begin
          $fwrite(f, "Register (34,15) Value: %h\n", PRED34_15_buffer[clk]);
        end
        if (PRED34_16_buffer[clk] != PRED34_16_buffer[!clk]) begin
          $fwrite(f, "Register (34,16) Value: %h\n", PRED34_16_buffer[clk]);
        end
        if (PRED34_17_buffer[clk] != PRED34_17_buffer[!clk]) begin
          $fwrite(f, "Register (34,17) Value: %h\n", PRED34_17_buffer[clk]);
        end
        if (PRED34_18_buffer[clk] != PRED34_18_buffer[!clk]) begin
          $fwrite(f, "Register (34,18) Value: %h\n", PRED34_18_buffer[clk]);
        end
        if (PRED34_19_buffer[clk] != PRED34_19_buffer[!clk]) begin
          $fwrite(f, "Register (34,19) Value: %h\n", PRED34_19_buffer[clk]);
        end
        if (PRED34_20_buffer[clk] != PRED34_20_buffer[!clk]) begin
          $fwrite(f, "Register (34,20) Value: %h\n", PRED34_20_buffer[clk]);
        end
        if (PRED34_21_buffer[clk] != PRED34_21_buffer[!clk]) begin
          $fwrite(f, "Register (34,21) Value: %h\n", PRED34_21_buffer[clk]);
        end
        if (PRED34_22_buffer[clk] != PRED34_22_buffer[!clk]) begin
          $fwrite(f, "Register (34,22) Value: %h\n", PRED34_22_buffer[clk]);
        end
        if (PRED34_23_buffer[clk] != PRED34_23_buffer[!clk]) begin
          $fwrite(f, "Register (34,23) Value: %h\n", PRED34_23_buffer[clk]);
        end
        if (PRED34_24_buffer[clk] != PRED34_24_buffer[!clk]) begin
          $fwrite(f, "Register (34,24) Value: %h\n", PRED34_24_buffer[clk]);
        end
        if (PRED34_25_buffer[clk] != PRED34_25_buffer[!clk]) begin
          $fwrite(f, "Register (34,25) Value: %h\n", PRED34_25_buffer[clk]);
        end
        if (PRED34_26_buffer[clk] != PRED34_26_buffer[!clk]) begin
          $fwrite(f, "Register (34,26) Value: %h\n", PRED34_26_buffer[clk]);
        end
        if (PRED34_27_buffer[clk] != PRED34_27_buffer[!clk]) begin
          $fwrite(f, "Register (34,27) Value: %h\n", PRED34_27_buffer[clk]);
        end
        if (PRED34_28_buffer[clk] != PRED34_28_buffer[!clk]) begin
          $fwrite(f, "Register (34,28) Value: %h\n", PRED34_28_buffer[clk]);
        end
        if (PRED34_29_buffer[clk] != PRED34_29_buffer[!clk]) begin
          $fwrite(f, "Register (34,29) Value: %h\n", PRED34_29_buffer[clk]);
        end
        if (PRED34_30_buffer[clk] != PRED34_30_buffer[!clk]) begin
          $fwrite(f, "Register (34,30) Value: %h\n", PRED34_30_buffer[clk]);
        end
        if (PRED34_31_buffer[clk] != PRED34_31_buffer[!clk]) begin
          $fwrite(f, "Register (34,31) Value: %h\n", PRED34_31_buffer[clk]);
        end
        if (PRED35_0_buffer[clk] != PRED35_0_buffer[!clk]) begin
          $fwrite(f, "Register (35,0) Value: %h\n", PRED35_0_buffer[clk]);
        end
        if (PRED35_1_buffer[clk] != PRED35_1_buffer[!clk]) begin
          $fwrite(f, "Register (35,1) Value: %h\n", PRED35_1_buffer[clk]);
        end
        if (PRED35_2_buffer[clk] != PRED35_2_buffer[!clk]) begin
          $fwrite(f, "Register (35,2) Value: %h\n", PRED35_2_buffer[clk]);
        end
        if (PRED35_3_buffer[clk] != PRED35_3_buffer[!clk]) begin
          $fwrite(f, "Register (35,3) Value: %h\n", PRED35_3_buffer[clk]);
        end
        if (PRED35_4_buffer[clk] != PRED35_4_buffer[!clk]) begin
          $fwrite(f, "Register (35,4) Value: %h\n", PRED35_4_buffer[clk]);
        end
        if (PRED35_5_buffer[clk] != PRED35_5_buffer[!clk]) begin
          $fwrite(f, "Register (35,5) Value: %h\n", PRED35_5_buffer[clk]);
        end
        if (PRED35_6_buffer[clk] != PRED35_6_buffer[!clk]) begin
          $fwrite(f, "Register (35,6) Value: %h\n", PRED35_6_buffer[clk]);
        end
        if (PRED35_7_buffer[clk] != PRED35_7_buffer[!clk]) begin
          $fwrite(f, "Register (35,7) Value: %h\n", PRED35_7_buffer[clk]);
        end
        if (PRED35_8_buffer[clk] != PRED35_8_buffer[!clk]) begin
          $fwrite(f, "Register (35,8) Value: %h\n", PRED35_8_buffer[clk]);
        end
        if (PRED35_9_buffer[clk] != PRED35_9_buffer[!clk]) begin
          $fwrite(f, "Register (35,9) Value: %h\n", PRED35_9_buffer[clk]);
        end
        if (PRED35_10_buffer[clk] != PRED35_10_buffer[!clk]) begin
          $fwrite(f, "Register (35,10) Value: %h\n", PRED35_10_buffer[clk]);
        end
        if (PRED35_11_buffer[clk] != PRED35_11_buffer[!clk]) begin
          $fwrite(f, "Register (35,11) Value: %h\n", PRED35_11_buffer[clk]);
        end
        if (PRED35_12_buffer[clk] != PRED35_12_buffer[!clk]) begin
          $fwrite(f, "Register (35,12) Value: %h\n", PRED35_12_buffer[clk]);
        end
        if (PRED35_13_buffer[clk] != PRED35_13_buffer[!clk]) begin
          $fwrite(f, "Register (35,13) Value: %h\n", PRED35_13_buffer[clk]);
        end
        if (PRED35_14_buffer[clk] != PRED35_14_buffer[!clk]) begin
          $fwrite(f, "Register (35,14) Value: %h\n", PRED35_14_buffer[clk]);
        end
        if (PRED35_15_buffer[clk] != PRED35_15_buffer[!clk]) begin
          $fwrite(f, "Register (35,15) Value: %h\n", PRED35_15_buffer[clk]);
        end
        if (PRED35_16_buffer[clk] != PRED35_16_buffer[!clk]) begin
          $fwrite(f, "Register (35,16) Value: %h\n", PRED35_16_buffer[clk]);
        end
        if (PRED35_17_buffer[clk] != PRED35_17_buffer[!clk]) begin
          $fwrite(f, "Register (35,17) Value: %h\n", PRED35_17_buffer[clk]);
        end
        if (PRED35_18_buffer[clk] != PRED35_18_buffer[!clk]) begin
          $fwrite(f, "Register (35,18) Value: %h\n", PRED35_18_buffer[clk]);
        end
        if (PRED35_19_buffer[clk] != PRED35_19_buffer[!clk]) begin
          $fwrite(f, "Register (35,19) Value: %h\n", PRED35_19_buffer[clk]);
        end
        if (PRED35_20_buffer[clk] != PRED35_20_buffer[!clk]) begin
          $fwrite(f, "Register (35,20) Value: %h\n", PRED35_20_buffer[clk]);
        end
        if (PRED35_21_buffer[clk] != PRED35_21_buffer[!clk]) begin
          $fwrite(f, "Register (35,21) Value: %h\n", PRED35_21_buffer[clk]);
        end
        if (PRED35_22_buffer[clk] != PRED35_22_buffer[!clk]) begin
          $fwrite(f, "Register (35,22) Value: %h\n", PRED35_22_buffer[clk]);
        end
        if (PRED35_23_buffer[clk] != PRED35_23_buffer[!clk]) begin
          $fwrite(f, "Register (35,23) Value: %h\n", PRED35_23_buffer[clk]);
        end
        if (PRED35_24_buffer[clk] != PRED35_24_buffer[!clk]) begin
          $fwrite(f, "Register (35,24) Value: %h\n", PRED35_24_buffer[clk]);
        end
        if (PRED35_25_buffer[clk] != PRED35_25_buffer[!clk]) begin
          $fwrite(f, "Register (35,25) Value: %h\n", PRED35_25_buffer[clk]);
        end
        if (PRED35_26_buffer[clk] != PRED35_26_buffer[!clk]) begin
          $fwrite(f, "Register (35,26) Value: %h\n", PRED35_26_buffer[clk]);
        end
        if (PRED35_27_buffer[clk] != PRED35_27_buffer[!clk]) begin
          $fwrite(f, "Register (35,27) Value: %h\n", PRED35_27_buffer[clk]);
        end
        if (PRED35_28_buffer[clk] != PRED35_28_buffer[!clk]) begin
          $fwrite(f, "Register (35,28) Value: %h\n", PRED35_28_buffer[clk]);
        end
        if (PRED35_29_buffer[clk] != PRED35_29_buffer[!clk]) begin
          $fwrite(f, "Register (35,29) Value: %h\n", PRED35_29_buffer[clk]);
        end
        if (PRED35_30_buffer[clk] != PRED35_30_buffer[!clk]) begin
          $fwrite(f, "Register (35,30) Value: %h\n", PRED35_30_buffer[clk]);
        end
        if (PRED35_31_buffer[clk] != PRED35_31_buffer[!clk]) begin
          $fwrite(f, "Register (35,31) Value: %h\n", PRED35_31_buffer[clk]);
        end
        if (PRED36_0_buffer[clk] != PRED36_0_buffer[!clk]) begin
          $fwrite(f, "Register (36,0) Value: %h\n", PRED36_0_buffer[clk]);
        end
        if (PRED36_1_buffer[clk] != PRED36_1_buffer[!clk]) begin
          $fwrite(f, "Register (36,1) Value: %h\n", PRED36_1_buffer[clk]);
        end
        if (PRED36_2_buffer[clk] != PRED36_2_buffer[!clk]) begin
          $fwrite(f, "Register (36,2) Value: %h\n", PRED36_2_buffer[clk]);
        end
        if (PRED36_3_buffer[clk] != PRED36_3_buffer[!clk]) begin
          $fwrite(f, "Register (36,3) Value: %h\n", PRED36_3_buffer[clk]);
        end
        if (PRED36_4_buffer[clk] != PRED36_4_buffer[!clk]) begin
          $fwrite(f, "Register (36,4) Value: %h\n", PRED36_4_buffer[clk]);
        end
        if (PRED36_5_buffer[clk] != PRED36_5_buffer[!clk]) begin
          $fwrite(f, "Register (36,5) Value: %h\n", PRED36_5_buffer[clk]);
        end
        if (PRED36_6_buffer[clk] != PRED36_6_buffer[!clk]) begin
          $fwrite(f, "Register (36,6) Value: %h\n", PRED36_6_buffer[clk]);
        end
        if (PRED36_7_buffer[clk] != PRED36_7_buffer[!clk]) begin
          $fwrite(f, "Register (36,7) Value: %h\n", PRED36_7_buffer[clk]);
        end
        if (PRED36_8_buffer[clk] != PRED36_8_buffer[!clk]) begin
          $fwrite(f, "Register (36,8) Value: %h\n", PRED36_8_buffer[clk]);
        end
        if (PRED36_9_buffer[clk] != PRED36_9_buffer[!clk]) begin
          $fwrite(f, "Register (36,9) Value: %h\n", PRED36_9_buffer[clk]);
        end
        if (PRED36_10_buffer[clk] != PRED36_10_buffer[!clk]) begin
          $fwrite(f, "Register (36,10) Value: %h\n", PRED36_10_buffer[clk]);
        end
        if (PRED36_11_buffer[clk] != PRED36_11_buffer[!clk]) begin
          $fwrite(f, "Register (36,11) Value: %h\n", PRED36_11_buffer[clk]);
        end
        if (PRED36_12_buffer[clk] != PRED36_12_buffer[!clk]) begin
          $fwrite(f, "Register (36,12) Value: %h\n", PRED36_12_buffer[clk]);
        end
        if (PRED36_13_buffer[clk] != PRED36_13_buffer[!clk]) begin
          $fwrite(f, "Register (36,13) Value: %h\n", PRED36_13_buffer[clk]);
        end
        if (PRED36_14_buffer[clk] != PRED36_14_buffer[!clk]) begin
          $fwrite(f, "Register (36,14) Value: %h\n", PRED36_14_buffer[clk]);
        end
        if (PRED36_15_buffer[clk] != PRED36_15_buffer[!clk]) begin
          $fwrite(f, "Register (36,15) Value: %h\n", PRED36_15_buffer[clk]);
        end
        if (PRED36_16_buffer[clk] != PRED36_16_buffer[!clk]) begin
          $fwrite(f, "Register (36,16) Value: %h\n", PRED36_16_buffer[clk]);
        end
        if (PRED36_17_buffer[clk] != PRED36_17_buffer[!clk]) begin
          $fwrite(f, "Register (36,17) Value: %h\n", PRED36_17_buffer[clk]);
        end
        if (PRED36_18_buffer[clk] != PRED36_18_buffer[!clk]) begin
          $fwrite(f, "Register (36,18) Value: %h\n", PRED36_18_buffer[clk]);
        end
        if (PRED36_19_buffer[clk] != PRED36_19_buffer[!clk]) begin
          $fwrite(f, "Register (36,19) Value: %h\n", PRED36_19_buffer[clk]);
        end
        if (PRED36_20_buffer[clk] != PRED36_20_buffer[!clk]) begin
          $fwrite(f, "Register (36,20) Value: %h\n", PRED36_20_buffer[clk]);
        end
        if (PRED36_21_buffer[clk] != PRED36_21_buffer[!clk]) begin
          $fwrite(f, "Register (36,21) Value: %h\n", PRED36_21_buffer[clk]);
        end
        if (PRED36_22_buffer[clk] != PRED36_22_buffer[!clk]) begin
          $fwrite(f, "Register (36,22) Value: %h\n", PRED36_22_buffer[clk]);
        end
        if (PRED36_23_buffer[clk] != PRED36_23_buffer[!clk]) begin
          $fwrite(f, "Register (36,23) Value: %h\n", PRED36_23_buffer[clk]);
        end
        if (PRED36_24_buffer[clk] != PRED36_24_buffer[!clk]) begin
          $fwrite(f, "Register (36,24) Value: %h\n", PRED36_24_buffer[clk]);
        end
        if (PRED36_25_buffer[clk] != PRED36_25_buffer[!clk]) begin
          $fwrite(f, "Register (36,25) Value: %h\n", PRED36_25_buffer[clk]);
        end
        if (PRED36_26_buffer[clk] != PRED36_26_buffer[!clk]) begin
          $fwrite(f, "Register (36,26) Value: %h\n", PRED36_26_buffer[clk]);
        end
        if (PRED36_27_buffer[clk] != PRED36_27_buffer[!clk]) begin
          $fwrite(f, "Register (36,27) Value: %h\n", PRED36_27_buffer[clk]);
        end
        if (PRED36_28_buffer[clk] != PRED36_28_buffer[!clk]) begin
          $fwrite(f, "Register (36,28) Value: %h\n", PRED36_28_buffer[clk]);
        end
        if (PRED36_29_buffer[clk] != PRED36_29_buffer[!clk]) begin
          $fwrite(f, "Register (36,29) Value: %h\n", PRED36_29_buffer[clk]);
        end
        if (PRED36_30_buffer[clk] != PRED36_30_buffer[!clk]) begin
          $fwrite(f, "Register (36,30) Value: %h\n", PRED36_30_buffer[clk]);
        end
        if (PRED36_31_buffer[clk] != PRED36_31_buffer[!clk]) begin
          $fwrite(f, "Register (36,31) Value: %h\n", PRED36_31_buffer[clk]);
        end
        if (PRED37_0_buffer[clk] != PRED37_0_buffer[!clk]) begin
          $fwrite(f, "Register (37,0) Value: %h\n", PRED37_0_buffer[clk]);
        end
        if (PRED37_1_buffer[clk] != PRED37_1_buffer[!clk]) begin
          $fwrite(f, "Register (37,1) Value: %h\n", PRED37_1_buffer[clk]);
        end
        if (PRED37_2_buffer[clk] != PRED37_2_buffer[!clk]) begin
          $fwrite(f, "Register (37,2) Value: %h\n", PRED37_2_buffer[clk]);
        end
        if (PRED37_3_buffer[clk] != PRED37_3_buffer[!clk]) begin
          $fwrite(f, "Register (37,3) Value: %h\n", PRED37_3_buffer[clk]);
        end
        if (PRED37_4_buffer[clk] != PRED37_4_buffer[!clk]) begin
          $fwrite(f, "Register (37,4) Value: %h\n", PRED37_4_buffer[clk]);
        end
        if (PRED37_5_buffer[clk] != PRED37_5_buffer[!clk]) begin
          $fwrite(f, "Register (37,5) Value: %h\n", PRED37_5_buffer[clk]);
        end
        if (PRED37_6_buffer[clk] != PRED37_6_buffer[!clk]) begin
          $fwrite(f, "Register (37,6) Value: %h\n", PRED37_6_buffer[clk]);
        end
        if (PRED37_7_buffer[clk] != PRED37_7_buffer[!clk]) begin
          $fwrite(f, "Register (37,7) Value: %h\n", PRED37_7_buffer[clk]);
        end
        if (PRED37_8_buffer[clk] != PRED37_8_buffer[!clk]) begin
          $fwrite(f, "Register (37,8) Value: %h\n", PRED37_8_buffer[clk]);
        end
        if (PRED37_9_buffer[clk] != PRED37_9_buffer[!clk]) begin
          $fwrite(f, "Register (37,9) Value: %h\n", PRED37_9_buffer[clk]);
        end
        if (PRED37_10_buffer[clk] != PRED37_10_buffer[!clk]) begin
          $fwrite(f, "Register (37,10) Value: %h\n", PRED37_10_buffer[clk]);
        end
        if (PRED37_11_buffer[clk] != PRED37_11_buffer[!clk]) begin
          $fwrite(f, "Register (37,11) Value: %h\n", PRED37_11_buffer[clk]);
        end
        if (PRED37_12_buffer[clk] != PRED37_12_buffer[!clk]) begin
          $fwrite(f, "Register (37,12) Value: %h\n", PRED37_12_buffer[clk]);
        end
        if (PRED37_13_buffer[clk] != PRED37_13_buffer[!clk]) begin
          $fwrite(f, "Register (37,13) Value: %h\n", PRED37_13_buffer[clk]);
        end
        if (PRED37_14_buffer[clk] != PRED37_14_buffer[!clk]) begin
          $fwrite(f, "Register (37,14) Value: %h\n", PRED37_14_buffer[clk]);
        end
        if (PRED37_15_buffer[clk] != PRED37_15_buffer[!clk]) begin
          $fwrite(f, "Register (37,15) Value: %h\n", PRED37_15_buffer[clk]);
        end
        if (PRED37_16_buffer[clk] != PRED37_16_buffer[!clk]) begin
          $fwrite(f, "Register (37,16) Value: %h\n", PRED37_16_buffer[clk]);
        end
        if (PRED37_17_buffer[clk] != PRED37_17_buffer[!clk]) begin
          $fwrite(f, "Register (37,17) Value: %h\n", PRED37_17_buffer[clk]);
        end
        if (PRED37_18_buffer[clk] != PRED37_18_buffer[!clk]) begin
          $fwrite(f, "Register (37,18) Value: %h\n", PRED37_18_buffer[clk]);
        end
        if (PRED37_19_buffer[clk] != PRED37_19_buffer[!clk]) begin
          $fwrite(f, "Register (37,19) Value: %h\n", PRED37_19_buffer[clk]);
        end
        if (PRED37_20_buffer[clk] != PRED37_20_buffer[!clk]) begin
          $fwrite(f, "Register (37,20) Value: %h\n", PRED37_20_buffer[clk]);
        end
        if (PRED37_21_buffer[clk] != PRED37_21_buffer[!clk]) begin
          $fwrite(f, "Register (37,21) Value: %h\n", PRED37_21_buffer[clk]);
        end
        if (PRED37_22_buffer[clk] != PRED37_22_buffer[!clk]) begin
          $fwrite(f, "Register (37,22) Value: %h\n", PRED37_22_buffer[clk]);
        end
        if (PRED37_23_buffer[clk] != PRED37_23_buffer[!clk]) begin
          $fwrite(f, "Register (37,23) Value: %h\n", PRED37_23_buffer[clk]);
        end
        if (PRED37_24_buffer[clk] != PRED37_24_buffer[!clk]) begin
          $fwrite(f, "Register (37,24) Value: %h\n", PRED37_24_buffer[clk]);
        end
        if (PRED37_25_buffer[clk] != PRED37_25_buffer[!clk]) begin
          $fwrite(f, "Register (37,25) Value: %h\n", PRED37_25_buffer[clk]);
        end
        if (PRED37_26_buffer[clk] != PRED37_26_buffer[!clk]) begin
          $fwrite(f, "Register (37,26) Value: %h\n", PRED37_26_buffer[clk]);
        end
        if (PRED37_27_buffer[clk] != PRED37_27_buffer[!clk]) begin
          $fwrite(f, "Register (37,27) Value: %h\n", PRED37_27_buffer[clk]);
        end
        if (PRED37_28_buffer[clk] != PRED37_28_buffer[!clk]) begin
          $fwrite(f, "Register (37,28) Value: %h\n", PRED37_28_buffer[clk]);
        end
        if (PRED37_29_buffer[clk] != PRED37_29_buffer[!clk]) begin
          $fwrite(f, "Register (37,29) Value: %h\n", PRED37_29_buffer[clk]);
        end
        if (PRED37_30_buffer[clk] != PRED37_30_buffer[!clk]) begin
          $fwrite(f, "Register (37,30) Value: %h\n", PRED37_30_buffer[clk]);
        end
        if (PRED37_31_buffer[clk] != PRED37_31_buffer[!clk]) begin
          $fwrite(f, "Register (37,31) Value: %h\n", PRED37_31_buffer[clk]);
        end
        if (PRED38_0_buffer[clk] != PRED38_0_buffer[!clk]) begin
          $fwrite(f, "Register (38,0) Value: %h\n", PRED38_0_buffer[clk]);
        end
        if (PRED38_1_buffer[clk] != PRED38_1_buffer[!clk]) begin
          $fwrite(f, "Register (38,1) Value: %h\n", PRED38_1_buffer[clk]);
        end
        if (PRED38_2_buffer[clk] != PRED38_2_buffer[!clk]) begin
          $fwrite(f, "Register (38,2) Value: %h\n", PRED38_2_buffer[clk]);
        end
        if (PRED38_3_buffer[clk] != PRED38_3_buffer[!clk]) begin
          $fwrite(f, "Register (38,3) Value: %h\n", PRED38_3_buffer[clk]);
        end
        if (PRED38_4_buffer[clk] != PRED38_4_buffer[!clk]) begin
          $fwrite(f, "Register (38,4) Value: %h\n", PRED38_4_buffer[clk]);
        end
        if (PRED38_5_buffer[clk] != PRED38_5_buffer[!clk]) begin
          $fwrite(f, "Register (38,5) Value: %h\n", PRED38_5_buffer[clk]);
        end
        if (PRED38_6_buffer[clk] != PRED38_6_buffer[!clk]) begin
          $fwrite(f, "Register (38,6) Value: %h\n", PRED38_6_buffer[clk]);
        end
        if (PRED38_7_buffer[clk] != PRED38_7_buffer[!clk]) begin
          $fwrite(f, "Register (38,7) Value: %h\n", PRED38_7_buffer[clk]);
        end
        if (PRED38_8_buffer[clk] != PRED38_8_buffer[!clk]) begin
          $fwrite(f, "Register (38,8) Value: %h\n", PRED38_8_buffer[clk]);
        end
        if (PRED38_9_buffer[clk] != PRED38_9_buffer[!clk]) begin
          $fwrite(f, "Register (38,9) Value: %h\n", PRED38_9_buffer[clk]);
        end
        if (PRED38_10_buffer[clk] != PRED38_10_buffer[!clk]) begin
          $fwrite(f, "Register (38,10) Value: %h\n", PRED38_10_buffer[clk]);
        end
        if (PRED38_11_buffer[clk] != PRED38_11_buffer[!clk]) begin
          $fwrite(f, "Register (38,11) Value: %h\n", PRED38_11_buffer[clk]);
        end
        if (PRED38_12_buffer[clk] != PRED38_12_buffer[!clk]) begin
          $fwrite(f, "Register (38,12) Value: %h\n", PRED38_12_buffer[clk]);
        end
        if (PRED38_13_buffer[clk] != PRED38_13_buffer[!clk]) begin
          $fwrite(f, "Register (38,13) Value: %h\n", PRED38_13_buffer[clk]);
        end
        if (PRED38_14_buffer[clk] != PRED38_14_buffer[!clk]) begin
          $fwrite(f, "Register (38,14) Value: %h\n", PRED38_14_buffer[clk]);
        end
        if (PRED38_15_buffer[clk] != PRED38_15_buffer[!clk]) begin
          $fwrite(f, "Register (38,15) Value: %h\n", PRED38_15_buffer[clk]);
        end
        if (PRED38_16_buffer[clk] != PRED38_16_buffer[!clk]) begin
          $fwrite(f, "Register (38,16) Value: %h\n", PRED38_16_buffer[clk]);
        end
        if (PRED38_17_buffer[clk] != PRED38_17_buffer[!clk]) begin
          $fwrite(f, "Register (38,17) Value: %h\n", PRED38_17_buffer[clk]);
        end
        if (PRED38_18_buffer[clk] != PRED38_18_buffer[!clk]) begin
          $fwrite(f, "Register (38,18) Value: %h\n", PRED38_18_buffer[clk]);
        end
        if (PRED38_19_buffer[clk] != PRED38_19_buffer[!clk]) begin
          $fwrite(f, "Register (38,19) Value: %h\n", PRED38_19_buffer[clk]);
        end
        if (PRED38_20_buffer[clk] != PRED38_20_buffer[!clk]) begin
          $fwrite(f, "Register (38,20) Value: %h\n", PRED38_20_buffer[clk]);
        end
        if (PRED38_21_buffer[clk] != PRED38_21_buffer[!clk]) begin
          $fwrite(f, "Register (38,21) Value: %h\n", PRED38_21_buffer[clk]);
        end
        if (PRED38_22_buffer[clk] != PRED38_22_buffer[!clk]) begin
          $fwrite(f, "Register (38,22) Value: %h\n", PRED38_22_buffer[clk]);
        end
        if (PRED38_23_buffer[clk] != PRED38_23_buffer[!clk]) begin
          $fwrite(f, "Register (38,23) Value: %h\n", PRED38_23_buffer[clk]);
        end
        if (PRED38_24_buffer[clk] != PRED38_24_buffer[!clk]) begin
          $fwrite(f, "Register (38,24) Value: %h\n", PRED38_24_buffer[clk]);
        end
        if (PRED38_25_buffer[clk] != PRED38_25_buffer[!clk]) begin
          $fwrite(f, "Register (38,25) Value: %h\n", PRED38_25_buffer[clk]);
        end
        if (PRED38_26_buffer[clk] != PRED38_26_buffer[!clk]) begin
          $fwrite(f, "Register (38,26) Value: %h\n", PRED38_26_buffer[clk]);
        end
        if (PRED38_27_buffer[clk] != PRED38_27_buffer[!clk]) begin
          $fwrite(f, "Register (38,27) Value: %h\n", PRED38_27_buffer[clk]);
        end
        if (PRED38_28_buffer[clk] != PRED38_28_buffer[!clk]) begin
          $fwrite(f, "Register (38,28) Value: %h\n", PRED38_28_buffer[clk]);
        end
        if (PRED38_29_buffer[clk] != PRED38_29_buffer[!clk]) begin
          $fwrite(f, "Register (38,29) Value: %h\n", PRED38_29_buffer[clk]);
        end
        if (PRED38_30_buffer[clk] != PRED38_30_buffer[!clk]) begin
          $fwrite(f, "Register (38,30) Value: %h\n", PRED38_30_buffer[clk]);
        end
        if (PRED38_31_buffer[clk] != PRED38_31_buffer[!clk]) begin
          $fwrite(f, "Register (38,31) Value: %h\n", PRED38_31_buffer[clk]);
        end
        if (PRED39_0_buffer[clk] != PRED39_0_buffer[!clk]) begin
          $fwrite(f, "Register (39,0) Value: %h\n", PRED39_0_buffer[clk]);
        end
        if (PRED39_1_buffer[clk] != PRED39_1_buffer[!clk]) begin
          $fwrite(f, "Register (39,1) Value: %h\n", PRED39_1_buffer[clk]);
        end
        if (PRED39_2_buffer[clk] != PRED39_2_buffer[!clk]) begin
          $fwrite(f, "Register (39,2) Value: %h\n", PRED39_2_buffer[clk]);
        end
        if (PRED39_3_buffer[clk] != PRED39_3_buffer[!clk]) begin
          $fwrite(f, "Register (39,3) Value: %h\n", PRED39_3_buffer[clk]);
        end
        if (PRED39_4_buffer[clk] != PRED39_4_buffer[!clk]) begin
          $fwrite(f, "Register (39,4) Value: %h\n", PRED39_4_buffer[clk]);
        end
        if (PRED39_5_buffer[clk] != PRED39_5_buffer[!clk]) begin
          $fwrite(f, "Register (39,5) Value: %h\n", PRED39_5_buffer[clk]);
        end
        if (PRED39_6_buffer[clk] != PRED39_6_buffer[!clk]) begin
          $fwrite(f, "Register (39,6) Value: %h\n", PRED39_6_buffer[clk]);
        end
        if (PRED39_7_buffer[clk] != PRED39_7_buffer[!clk]) begin
          $fwrite(f, "Register (39,7) Value: %h\n", PRED39_7_buffer[clk]);
        end
        if (PRED39_8_buffer[clk] != PRED39_8_buffer[!clk]) begin
          $fwrite(f, "Register (39,8) Value: %h\n", PRED39_8_buffer[clk]);
        end
        if (PRED39_9_buffer[clk] != PRED39_9_buffer[!clk]) begin
          $fwrite(f, "Register (39,9) Value: %h\n", PRED39_9_buffer[clk]);
        end
        if (PRED39_10_buffer[clk] != PRED39_10_buffer[!clk]) begin
          $fwrite(f, "Register (39,10) Value: %h\n", PRED39_10_buffer[clk]);
        end
        if (PRED39_11_buffer[clk] != PRED39_11_buffer[!clk]) begin
          $fwrite(f, "Register (39,11) Value: %h\n", PRED39_11_buffer[clk]);
        end
        if (PRED39_12_buffer[clk] != PRED39_12_buffer[!clk]) begin
          $fwrite(f, "Register (39,12) Value: %h\n", PRED39_12_buffer[clk]);
        end
        if (PRED39_13_buffer[clk] != PRED39_13_buffer[!clk]) begin
          $fwrite(f, "Register (39,13) Value: %h\n", PRED39_13_buffer[clk]);
        end
        if (PRED39_14_buffer[clk] != PRED39_14_buffer[!clk]) begin
          $fwrite(f, "Register (39,14) Value: %h\n", PRED39_14_buffer[clk]);
        end
        if (PRED39_15_buffer[clk] != PRED39_15_buffer[!clk]) begin
          $fwrite(f, "Register (39,15) Value: %h\n", PRED39_15_buffer[clk]);
        end
        if (PRED39_16_buffer[clk] != PRED39_16_buffer[!clk]) begin
          $fwrite(f, "Register (39,16) Value: %h\n", PRED39_16_buffer[clk]);
        end
        if (PRED39_17_buffer[clk] != PRED39_17_buffer[!clk]) begin
          $fwrite(f, "Register (39,17) Value: %h\n", PRED39_17_buffer[clk]);
        end
        if (PRED39_18_buffer[clk] != PRED39_18_buffer[!clk]) begin
          $fwrite(f, "Register (39,18) Value: %h\n", PRED39_18_buffer[clk]);
        end
        if (PRED39_19_buffer[clk] != PRED39_19_buffer[!clk]) begin
          $fwrite(f, "Register (39,19) Value: %h\n", PRED39_19_buffer[clk]);
        end
        if (PRED39_20_buffer[clk] != PRED39_20_buffer[!clk]) begin
          $fwrite(f, "Register (39,20) Value: %h\n", PRED39_20_buffer[clk]);
        end
        if (PRED39_21_buffer[clk] != PRED39_21_buffer[!clk]) begin
          $fwrite(f, "Register (39,21) Value: %h\n", PRED39_21_buffer[clk]);
        end
        if (PRED39_22_buffer[clk] != PRED39_22_buffer[!clk]) begin
          $fwrite(f, "Register (39,22) Value: %h\n", PRED39_22_buffer[clk]);
        end
        if (PRED39_23_buffer[clk] != PRED39_23_buffer[!clk]) begin
          $fwrite(f, "Register (39,23) Value: %h\n", PRED39_23_buffer[clk]);
        end
        if (PRED39_24_buffer[clk] != PRED39_24_buffer[!clk]) begin
          $fwrite(f, "Register (39,24) Value: %h\n", PRED39_24_buffer[clk]);
        end
        if (PRED39_25_buffer[clk] != PRED39_25_buffer[!clk]) begin
          $fwrite(f, "Register (39,25) Value: %h\n", PRED39_25_buffer[clk]);
        end
        if (PRED39_26_buffer[clk] != PRED39_26_buffer[!clk]) begin
          $fwrite(f, "Register (39,26) Value: %h\n", PRED39_26_buffer[clk]);
        end
        if (PRED39_27_buffer[clk] != PRED39_27_buffer[!clk]) begin
          $fwrite(f, "Register (39,27) Value: %h\n", PRED39_27_buffer[clk]);
        end
        if (PRED39_28_buffer[clk] != PRED39_28_buffer[!clk]) begin
          $fwrite(f, "Register (39,28) Value: %h\n", PRED39_28_buffer[clk]);
        end
        if (PRED39_29_buffer[clk] != PRED39_29_buffer[!clk]) begin
          $fwrite(f, "Register (39,29) Value: %h\n", PRED39_29_buffer[clk]);
        end
        if (PRED39_30_buffer[clk] != PRED39_30_buffer[!clk]) begin
          $fwrite(f, "Register (39,30) Value: %h\n", PRED39_30_buffer[clk]);
        end
        if (PRED39_31_buffer[clk] != PRED39_31_buffer[!clk]) begin
          $fwrite(f, "Register (39,31) Value: %h\n", PRED39_31_buffer[clk]);
        end
        if (PRED40_0_buffer[clk] != PRED40_0_buffer[!clk]) begin
          $fwrite(f, "Register (40,0) Value: %h\n", PRED40_0_buffer[clk]);
        end
        if (PRED40_1_buffer[clk] != PRED40_1_buffer[!clk]) begin
          $fwrite(f, "Register (40,1) Value: %h\n", PRED40_1_buffer[clk]);
        end
        if (PRED40_2_buffer[clk] != PRED40_2_buffer[!clk]) begin
          $fwrite(f, "Register (40,2) Value: %h\n", PRED40_2_buffer[clk]);
        end
        if (PRED40_3_buffer[clk] != PRED40_3_buffer[!clk]) begin
          $fwrite(f, "Register (40,3) Value: %h\n", PRED40_3_buffer[clk]);
        end
        if (PRED40_4_buffer[clk] != PRED40_4_buffer[!clk]) begin
          $fwrite(f, "Register (40,4) Value: %h\n", PRED40_4_buffer[clk]);
        end
        if (PRED40_5_buffer[clk] != PRED40_5_buffer[!clk]) begin
          $fwrite(f, "Register (40,5) Value: %h\n", PRED40_5_buffer[clk]);
        end
        if (PRED40_6_buffer[clk] != PRED40_6_buffer[!clk]) begin
          $fwrite(f, "Register (40,6) Value: %h\n", PRED40_6_buffer[clk]);
        end
        if (PRED40_7_buffer[clk] != PRED40_7_buffer[!clk]) begin
          $fwrite(f, "Register (40,7) Value: %h\n", PRED40_7_buffer[clk]);
        end
        if (PRED40_8_buffer[clk] != PRED40_8_buffer[!clk]) begin
          $fwrite(f, "Register (40,8) Value: %h\n", PRED40_8_buffer[clk]);
        end
        if (PRED40_9_buffer[clk] != PRED40_9_buffer[!clk]) begin
          $fwrite(f, "Register (40,9) Value: %h\n", PRED40_9_buffer[clk]);
        end
        if (PRED40_10_buffer[clk] != PRED40_10_buffer[!clk]) begin
          $fwrite(f, "Register (40,10) Value: %h\n", PRED40_10_buffer[clk]);
        end
        if (PRED40_11_buffer[clk] != PRED40_11_buffer[!clk]) begin
          $fwrite(f, "Register (40,11) Value: %h\n", PRED40_11_buffer[clk]);
        end
        if (PRED40_12_buffer[clk] != PRED40_12_buffer[!clk]) begin
          $fwrite(f, "Register (40,12) Value: %h\n", PRED40_12_buffer[clk]);
        end
        if (PRED40_13_buffer[clk] != PRED40_13_buffer[!clk]) begin
          $fwrite(f, "Register (40,13) Value: %h\n", PRED40_13_buffer[clk]);
        end
        if (PRED40_14_buffer[clk] != PRED40_14_buffer[!clk]) begin
          $fwrite(f, "Register (40,14) Value: %h\n", PRED40_14_buffer[clk]);
        end
        if (PRED40_15_buffer[clk] != PRED40_15_buffer[!clk]) begin
          $fwrite(f, "Register (40,15) Value: %h\n", PRED40_15_buffer[clk]);
        end
        if (PRED40_16_buffer[clk] != PRED40_16_buffer[!clk]) begin
          $fwrite(f, "Register (40,16) Value: %h\n", PRED40_16_buffer[clk]);
        end
        if (PRED40_17_buffer[clk] != PRED40_17_buffer[!clk]) begin
          $fwrite(f, "Register (40,17) Value: %h\n", PRED40_17_buffer[clk]);
        end
        if (PRED40_18_buffer[clk] != PRED40_18_buffer[!clk]) begin
          $fwrite(f, "Register (40,18) Value: %h\n", PRED40_18_buffer[clk]);
        end
        if (PRED40_19_buffer[clk] != PRED40_19_buffer[!clk]) begin
          $fwrite(f, "Register (40,19) Value: %h\n", PRED40_19_buffer[clk]);
        end
        if (PRED40_20_buffer[clk] != PRED40_20_buffer[!clk]) begin
          $fwrite(f, "Register (40,20) Value: %h\n", PRED40_20_buffer[clk]);
        end
        if (PRED40_21_buffer[clk] != PRED40_21_buffer[!clk]) begin
          $fwrite(f, "Register (40,21) Value: %h\n", PRED40_21_buffer[clk]);
        end
        if (PRED40_22_buffer[clk] != PRED40_22_buffer[!clk]) begin
          $fwrite(f, "Register (40,22) Value: %h\n", PRED40_22_buffer[clk]);
        end
        if (PRED40_23_buffer[clk] != PRED40_23_buffer[!clk]) begin
          $fwrite(f, "Register (40,23) Value: %h\n", PRED40_23_buffer[clk]);
        end
        if (PRED40_24_buffer[clk] != PRED40_24_buffer[!clk]) begin
          $fwrite(f, "Register (40,24) Value: %h\n", PRED40_24_buffer[clk]);
        end
        if (PRED40_25_buffer[clk] != PRED40_25_buffer[!clk]) begin
          $fwrite(f, "Register (40,25) Value: %h\n", PRED40_25_buffer[clk]);
        end
        if (PRED40_26_buffer[clk] != PRED40_26_buffer[!clk]) begin
          $fwrite(f, "Register (40,26) Value: %h\n", PRED40_26_buffer[clk]);
        end
        if (PRED40_27_buffer[clk] != PRED40_27_buffer[!clk]) begin
          $fwrite(f, "Register (40,27) Value: %h\n", PRED40_27_buffer[clk]);
        end
        if (PRED40_28_buffer[clk] != PRED40_28_buffer[!clk]) begin
          $fwrite(f, "Register (40,28) Value: %h\n", PRED40_28_buffer[clk]);
        end
        if (PRED40_29_buffer[clk] != PRED40_29_buffer[!clk]) begin
          $fwrite(f, "Register (40,29) Value: %h\n", PRED40_29_buffer[clk]);
        end
        if (PRED40_30_buffer[clk] != PRED40_30_buffer[!clk]) begin
          $fwrite(f, "Register (40,30) Value: %h\n", PRED40_30_buffer[clk]);
        end
        if (PRED40_31_buffer[clk] != PRED40_31_buffer[!clk]) begin
          $fwrite(f, "Register (40,31) Value: %h\n", PRED40_31_buffer[clk]);
        end
        if (PRED41_0_buffer[clk] != PRED41_0_buffer[!clk]) begin
          $fwrite(f, "Register (41,0) Value: %h\n", PRED41_0_buffer[clk]);
        end
        if (PRED41_1_buffer[clk] != PRED41_1_buffer[!clk]) begin
          $fwrite(f, "Register (41,1) Value: %h\n", PRED41_1_buffer[clk]);
        end
        if (PRED41_2_buffer[clk] != PRED41_2_buffer[!clk]) begin
          $fwrite(f, "Register (41,2) Value: %h\n", PRED41_2_buffer[clk]);
        end
        if (PRED41_3_buffer[clk] != PRED41_3_buffer[!clk]) begin
          $fwrite(f, "Register (41,3) Value: %h\n", PRED41_3_buffer[clk]);
        end
        if (PRED41_4_buffer[clk] != PRED41_4_buffer[!clk]) begin
          $fwrite(f, "Register (41,4) Value: %h\n", PRED41_4_buffer[clk]);
        end
        if (PRED41_5_buffer[clk] != PRED41_5_buffer[!clk]) begin
          $fwrite(f, "Register (41,5) Value: %h\n", PRED41_5_buffer[clk]);
        end
        if (PRED41_6_buffer[clk] != PRED41_6_buffer[!clk]) begin
          $fwrite(f, "Register (41,6) Value: %h\n", PRED41_6_buffer[clk]);
        end
        if (PRED41_7_buffer[clk] != PRED41_7_buffer[!clk]) begin
          $fwrite(f, "Register (41,7) Value: %h\n", PRED41_7_buffer[clk]);
        end
        if (PRED41_8_buffer[clk] != PRED41_8_buffer[!clk]) begin
          $fwrite(f, "Register (41,8) Value: %h\n", PRED41_8_buffer[clk]);
        end
        if (PRED41_9_buffer[clk] != PRED41_9_buffer[!clk]) begin
          $fwrite(f, "Register (41,9) Value: %h\n", PRED41_9_buffer[clk]);
        end
        if (PRED41_10_buffer[clk] != PRED41_10_buffer[!clk]) begin
          $fwrite(f, "Register (41,10) Value: %h\n", PRED41_10_buffer[clk]);
        end
        if (PRED41_11_buffer[clk] != PRED41_11_buffer[!clk]) begin
          $fwrite(f, "Register (41,11) Value: %h\n", PRED41_11_buffer[clk]);
        end
        if (PRED41_12_buffer[clk] != PRED41_12_buffer[!clk]) begin
          $fwrite(f, "Register (41,12) Value: %h\n", PRED41_12_buffer[clk]);
        end
        if (PRED41_13_buffer[clk] != PRED41_13_buffer[!clk]) begin
          $fwrite(f, "Register (41,13) Value: %h\n", PRED41_13_buffer[clk]);
        end
        if (PRED41_14_buffer[clk] != PRED41_14_buffer[!clk]) begin
          $fwrite(f, "Register (41,14) Value: %h\n", PRED41_14_buffer[clk]);
        end
        if (PRED41_15_buffer[clk] != PRED41_15_buffer[!clk]) begin
          $fwrite(f, "Register (41,15) Value: %h\n", PRED41_15_buffer[clk]);
        end
        if (PRED41_16_buffer[clk] != PRED41_16_buffer[!clk]) begin
          $fwrite(f, "Register (41,16) Value: %h\n", PRED41_16_buffer[clk]);
        end
        if (PRED41_17_buffer[clk] != PRED41_17_buffer[!clk]) begin
          $fwrite(f, "Register (41,17) Value: %h\n", PRED41_17_buffer[clk]);
        end
        if (PRED41_18_buffer[clk] != PRED41_18_buffer[!clk]) begin
          $fwrite(f, "Register (41,18) Value: %h\n", PRED41_18_buffer[clk]);
        end
        if (PRED41_19_buffer[clk] != PRED41_19_buffer[!clk]) begin
          $fwrite(f, "Register (41,19) Value: %h\n", PRED41_19_buffer[clk]);
        end
        if (PRED41_20_buffer[clk] != PRED41_20_buffer[!clk]) begin
          $fwrite(f, "Register (41,20) Value: %h\n", PRED41_20_buffer[clk]);
        end
        if (PRED41_21_buffer[clk] != PRED41_21_buffer[!clk]) begin
          $fwrite(f, "Register (41,21) Value: %h\n", PRED41_21_buffer[clk]);
        end
        if (PRED41_22_buffer[clk] != PRED41_22_buffer[!clk]) begin
          $fwrite(f, "Register (41,22) Value: %h\n", PRED41_22_buffer[clk]);
        end
        if (PRED41_23_buffer[clk] != PRED41_23_buffer[!clk]) begin
          $fwrite(f, "Register (41,23) Value: %h\n", PRED41_23_buffer[clk]);
        end
        if (PRED41_24_buffer[clk] != PRED41_24_buffer[!clk]) begin
          $fwrite(f, "Register (41,24) Value: %h\n", PRED41_24_buffer[clk]);
        end
        if (PRED41_25_buffer[clk] != PRED41_25_buffer[!clk]) begin
          $fwrite(f, "Register (41,25) Value: %h\n", PRED41_25_buffer[clk]);
        end
        if (PRED41_26_buffer[clk] != PRED41_26_buffer[!clk]) begin
          $fwrite(f, "Register (41,26) Value: %h\n", PRED41_26_buffer[clk]);
        end
        if (PRED41_27_buffer[clk] != PRED41_27_buffer[!clk]) begin
          $fwrite(f, "Register (41,27) Value: %h\n", PRED41_27_buffer[clk]);
        end
        if (PRED41_28_buffer[clk] != PRED41_28_buffer[!clk]) begin
          $fwrite(f, "Register (41,28) Value: %h\n", PRED41_28_buffer[clk]);
        end
        if (PRED41_29_buffer[clk] != PRED41_29_buffer[!clk]) begin
          $fwrite(f, "Register (41,29) Value: %h\n", PRED41_29_buffer[clk]);
        end
        if (PRED41_30_buffer[clk] != PRED41_30_buffer[!clk]) begin
          $fwrite(f, "Register (41,30) Value: %h\n", PRED41_30_buffer[clk]);
        end
        if (PRED41_31_buffer[clk] != PRED41_31_buffer[!clk]) begin
          $fwrite(f, "Register (41,31) Value: %h\n", PRED41_31_buffer[clk]);
        end
        if (PRED42_0_buffer[clk] != PRED42_0_buffer[!clk]) begin
          $fwrite(f, "Register (42,0) Value: %h\n", PRED42_0_buffer[clk]);
        end
        if (PRED42_1_buffer[clk] != PRED42_1_buffer[!clk]) begin
          $fwrite(f, "Register (42,1) Value: %h\n", PRED42_1_buffer[clk]);
        end
        if (PRED42_2_buffer[clk] != PRED42_2_buffer[!clk]) begin
          $fwrite(f, "Register (42,2) Value: %h\n", PRED42_2_buffer[clk]);
        end
        if (PRED42_3_buffer[clk] != PRED42_3_buffer[!clk]) begin
          $fwrite(f, "Register (42,3) Value: %h\n", PRED42_3_buffer[clk]);
        end
        if (PRED42_4_buffer[clk] != PRED42_4_buffer[!clk]) begin
          $fwrite(f, "Register (42,4) Value: %h\n", PRED42_4_buffer[clk]);
        end
        if (PRED42_5_buffer[clk] != PRED42_5_buffer[!clk]) begin
          $fwrite(f, "Register (42,5) Value: %h\n", PRED42_5_buffer[clk]);
        end
        if (PRED42_6_buffer[clk] != PRED42_6_buffer[!clk]) begin
          $fwrite(f, "Register (42,6) Value: %h\n", PRED42_6_buffer[clk]);
        end
        if (PRED42_7_buffer[clk] != PRED42_7_buffer[!clk]) begin
          $fwrite(f, "Register (42,7) Value: %h\n", PRED42_7_buffer[clk]);
        end
        if (PRED42_8_buffer[clk] != PRED42_8_buffer[!clk]) begin
          $fwrite(f, "Register (42,8) Value: %h\n", PRED42_8_buffer[clk]);
        end
        if (PRED42_9_buffer[clk] != PRED42_9_buffer[!clk]) begin
          $fwrite(f, "Register (42,9) Value: %h\n", PRED42_9_buffer[clk]);
        end
        if (PRED42_10_buffer[clk] != PRED42_10_buffer[!clk]) begin
          $fwrite(f, "Register (42,10) Value: %h\n", PRED42_10_buffer[clk]);
        end
        if (PRED42_11_buffer[clk] != PRED42_11_buffer[!clk]) begin
          $fwrite(f, "Register (42,11) Value: %h\n", PRED42_11_buffer[clk]);
        end
        if (PRED42_12_buffer[clk] != PRED42_12_buffer[!clk]) begin
          $fwrite(f, "Register (42,12) Value: %h\n", PRED42_12_buffer[clk]);
        end
        if (PRED42_13_buffer[clk] != PRED42_13_buffer[!clk]) begin
          $fwrite(f, "Register (42,13) Value: %h\n", PRED42_13_buffer[clk]);
        end
        if (PRED42_14_buffer[clk] != PRED42_14_buffer[!clk]) begin
          $fwrite(f, "Register (42,14) Value: %h\n", PRED42_14_buffer[clk]);
        end
        if (PRED42_15_buffer[clk] != PRED42_15_buffer[!clk]) begin
          $fwrite(f, "Register (42,15) Value: %h\n", PRED42_15_buffer[clk]);
        end
        if (PRED42_16_buffer[clk] != PRED42_16_buffer[!clk]) begin
          $fwrite(f, "Register (42,16) Value: %h\n", PRED42_16_buffer[clk]);
        end
        if (PRED42_17_buffer[clk] != PRED42_17_buffer[!clk]) begin
          $fwrite(f, "Register (42,17) Value: %h\n", PRED42_17_buffer[clk]);
        end
        if (PRED42_18_buffer[clk] != PRED42_18_buffer[!clk]) begin
          $fwrite(f, "Register (42,18) Value: %h\n", PRED42_18_buffer[clk]);
        end
        if (PRED42_19_buffer[clk] != PRED42_19_buffer[!clk]) begin
          $fwrite(f, "Register (42,19) Value: %h\n", PRED42_19_buffer[clk]);
        end
        if (PRED42_20_buffer[clk] != PRED42_20_buffer[!clk]) begin
          $fwrite(f, "Register (42,20) Value: %h\n", PRED42_20_buffer[clk]);
        end
        if (PRED42_21_buffer[clk] != PRED42_21_buffer[!clk]) begin
          $fwrite(f, "Register (42,21) Value: %h\n", PRED42_21_buffer[clk]);
        end
        if (PRED42_22_buffer[clk] != PRED42_22_buffer[!clk]) begin
          $fwrite(f, "Register (42,22) Value: %h\n", PRED42_22_buffer[clk]);
        end
        if (PRED42_23_buffer[clk] != PRED42_23_buffer[!clk]) begin
          $fwrite(f, "Register (42,23) Value: %h\n", PRED42_23_buffer[clk]);
        end
        if (PRED42_24_buffer[clk] != PRED42_24_buffer[!clk]) begin
          $fwrite(f, "Register (42,24) Value: %h\n", PRED42_24_buffer[clk]);
        end
        if (PRED42_25_buffer[clk] != PRED42_25_buffer[!clk]) begin
          $fwrite(f, "Register (42,25) Value: %h\n", PRED42_25_buffer[clk]);
        end
        if (PRED42_26_buffer[clk] != PRED42_26_buffer[!clk]) begin
          $fwrite(f, "Register (42,26) Value: %h\n", PRED42_26_buffer[clk]);
        end
        if (PRED42_27_buffer[clk] != PRED42_27_buffer[!clk]) begin
          $fwrite(f, "Register (42,27) Value: %h\n", PRED42_27_buffer[clk]);
        end
        if (PRED42_28_buffer[clk] != PRED42_28_buffer[!clk]) begin
          $fwrite(f, "Register (42,28) Value: %h\n", PRED42_28_buffer[clk]);
        end
        if (PRED42_29_buffer[clk] != PRED42_29_buffer[!clk]) begin
          $fwrite(f, "Register (42,29) Value: %h\n", PRED42_29_buffer[clk]);
        end
        if (PRED42_30_buffer[clk] != PRED42_30_buffer[!clk]) begin
          $fwrite(f, "Register (42,30) Value: %h\n", PRED42_30_buffer[clk]);
        end
        if (PRED42_31_buffer[clk] != PRED42_31_buffer[!clk]) begin
          $fwrite(f, "Register (42,31) Value: %h\n", PRED42_31_buffer[clk]);
        end
        if (PRED43_0_buffer[clk] != PRED43_0_buffer[!clk]) begin
          $fwrite(f, "Register (43,0) Value: %h\n", PRED43_0_buffer[clk]);
        end
        if (PRED43_1_buffer[clk] != PRED43_1_buffer[!clk]) begin
          $fwrite(f, "Register (43,1) Value: %h\n", PRED43_1_buffer[clk]);
        end
        if (PRED43_2_buffer[clk] != PRED43_2_buffer[!clk]) begin
          $fwrite(f, "Register (43,2) Value: %h\n", PRED43_2_buffer[clk]);
        end
        if (PRED43_3_buffer[clk] != PRED43_3_buffer[!clk]) begin
          $fwrite(f, "Register (43,3) Value: %h\n", PRED43_3_buffer[clk]);
        end
        if (PRED43_4_buffer[clk] != PRED43_4_buffer[!clk]) begin
          $fwrite(f, "Register (43,4) Value: %h\n", PRED43_4_buffer[clk]);
        end
        if (PRED43_5_buffer[clk] != PRED43_5_buffer[!clk]) begin
          $fwrite(f, "Register (43,5) Value: %h\n", PRED43_5_buffer[clk]);
        end
        if (PRED43_6_buffer[clk] != PRED43_6_buffer[!clk]) begin
          $fwrite(f, "Register (43,6) Value: %h\n", PRED43_6_buffer[clk]);
        end
        if (PRED43_7_buffer[clk] != PRED43_7_buffer[!clk]) begin
          $fwrite(f, "Register (43,7) Value: %h\n", PRED43_7_buffer[clk]);
        end
        if (PRED43_8_buffer[clk] != PRED43_8_buffer[!clk]) begin
          $fwrite(f, "Register (43,8) Value: %h\n", PRED43_8_buffer[clk]);
        end
        if (PRED43_9_buffer[clk] != PRED43_9_buffer[!clk]) begin
          $fwrite(f, "Register (43,9) Value: %h\n", PRED43_9_buffer[clk]);
        end
        if (PRED43_10_buffer[clk] != PRED43_10_buffer[!clk]) begin
          $fwrite(f, "Register (43,10) Value: %h\n", PRED43_10_buffer[clk]);
        end
        if (PRED43_11_buffer[clk] != PRED43_11_buffer[!clk]) begin
          $fwrite(f, "Register (43,11) Value: %h\n", PRED43_11_buffer[clk]);
        end
        if (PRED43_12_buffer[clk] != PRED43_12_buffer[!clk]) begin
          $fwrite(f, "Register (43,12) Value: %h\n", PRED43_12_buffer[clk]);
        end
        if (PRED43_13_buffer[clk] != PRED43_13_buffer[!clk]) begin
          $fwrite(f, "Register (43,13) Value: %h\n", PRED43_13_buffer[clk]);
        end
        if (PRED43_14_buffer[clk] != PRED43_14_buffer[!clk]) begin
          $fwrite(f, "Register (43,14) Value: %h\n", PRED43_14_buffer[clk]);
        end
        if (PRED43_15_buffer[clk] != PRED43_15_buffer[!clk]) begin
          $fwrite(f, "Register (43,15) Value: %h\n", PRED43_15_buffer[clk]);
        end
        if (PRED43_16_buffer[clk] != PRED43_16_buffer[!clk]) begin
          $fwrite(f, "Register (43,16) Value: %h\n", PRED43_16_buffer[clk]);
        end
        if (PRED43_17_buffer[clk] != PRED43_17_buffer[!clk]) begin
          $fwrite(f, "Register (43,17) Value: %h\n", PRED43_17_buffer[clk]);
        end
        if (PRED43_18_buffer[clk] != PRED43_18_buffer[!clk]) begin
          $fwrite(f, "Register (43,18) Value: %h\n", PRED43_18_buffer[clk]);
        end
        if (PRED43_19_buffer[clk] != PRED43_19_buffer[!clk]) begin
          $fwrite(f, "Register (43,19) Value: %h\n", PRED43_19_buffer[clk]);
        end
        if (PRED43_20_buffer[clk] != PRED43_20_buffer[!clk]) begin
          $fwrite(f, "Register (43,20) Value: %h\n", PRED43_20_buffer[clk]);
        end
        if (PRED43_21_buffer[clk] != PRED43_21_buffer[!clk]) begin
          $fwrite(f, "Register (43,21) Value: %h\n", PRED43_21_buffer[clk]);
        end
        if (PRED43_22_buffer[clk] != PRED43_22_buffer[!clk]) begin
          $fwrite(f, "Register (43,22) Value: %h\n", PRED43_22_buffer[clk]);
        end
        if (PRED43_23_buffer[clk] != PRED43_23_buffer[!clk]) begin
          $fwrite(f, "Register (43,23) Value: %h\n", PRED43_23_buffer[clk]);
        end
        if (PRED43_24_buffer[clk] != PRED43_24_buffer[!clk]) begin
          $fwrite(f, "Register (43,24) Value: %h\n", PRED43_24_buffer[clk]);
        end
        if (PRED43_25_buffer[clk] != PRED43_25_buffer[!clk]) begin
          $fwrite(f, "Register (43,25) Value: %h\n", PRED43_25_buffer[clk]);
        end
        if (PRED43_26_buffer[clk] != PRED43_26_buffer[!clk]) begin
          $fwrite(f, "Register (43,26) Value: %h\n", PRED43_26_buffer[clk]);
        end
        if (PRED43_27_buffer[clk] != PRED43_27_buffer[!clk]) begin
          $fwrite(f, "Register (43,27) Value: %h\n", PRED43_27_buffer[clk]);
        end
        if (PRED43_28_buffer[clk] != PRED43_28_buffer[!clk]) begin
          $fwrite(f, "Register (43,28) Value: %h\n", PRED43_28_buffer[clk]);
        end
        if (PRED43_29_buffer[clk] != PRED43_29_buffer[!clk]) begin
          $fwrite(f, "Register (43,29) Value: %h\n", PRED43_29_buffer[clk]);
        end
        if (PRED43_30_buffer[clk] != PRED43_30_buffer[!clk]) begin
          $fwrite(f, "Register (43,30) Value: %h\n", PRED43_30_buffer[clk]);
        end
        if (PRED43_31_buffer[clk] != PRED43_31_buffer[!clk]) begin
          $fwrite(f, "Register (43,31) Value: %h\n", PRED43_31_buffer[clk]);
        end
        if (PRED44_0_buffer[clk] != PRED44_0_buffer[!clk]) begin
          $fwrite(f, "Register (44,0) Value: %h\n", PRED44_0_buffer[clk]);
        end
        if (PRED44_1_buffer[clk] != PRED44_1_buffer[!clk]) begin
          $fwrite(f, "Register (44,1) Value: %h\n", PRED44_1_buffer[clk]);
        end
        if (PRED44_2_buffer[clk] != PRED44_2_buffer[!clk]) begin
          $fwrite(f, "Register (44,2) Value: %h\n", PRED44_2_buffer[clk]);
        end
        if (PRED44_3_buffer[clk] != PRED44_3_buffer[!clk]) begin
          $fwrite(f, "Register (44,3) Value: %h\n", PRED44_3_buffer[clk]);
        end
        if (PRED44_4_buffer[clk] != PRED44_4_buffer[!clk]) begin
          $fwrite(f, "Register (44,4) Value: %h\n", PRED44_4_buffer[clk]);
        end
        if (PRED44_5_buffer[clk] != PRED44_5_buffer[!clk]) begin
          $fwrite(f, "Register (44,5) Value: %h\n", PRED44_5_buffer[clk]);
        end
        if (PRED44_6_buffer[clk] != PRED44_6_buffer[!clk]) begin
          $fwrite(f, "Register (44,6) Value: %h\n", PRED44_6_buffer[clk]);
        end
        if (PRED44_7_buffer[clk] != PRED44_7_buffer[!clk]) begin
          $fwrite(f, "Register (44,7) Value: %h\n", PRED44_7_buffer[clk]);
        end
        if (PRED44_8_buffer[clk] != PRED44_8_buffer[!clk]) begin
          $fwrite(f, "Register (44,8) Value: %h\n", PRED44_8_buffer[clk]);
        end
        if (PRED44_9_buffer[clk] != PRED44_9_buffer[!clk]) begin
          $fwrite(f, "Register (44,9) Value: %h\n", PRED44_9_buffer[clk]);
        end
        if (PRED44_10_buffer[clk] != PRED44_10_buffer[!clk]) begin
          $fwrite(f, "Register (44,10) Value: %h\n", PRED44_10_buffer[clk]);
        end
        if (PRED44_11_buffer[clk] != PRED44_11_buffer[!clk]) begin
          $fwrite(f, "Register (44,11) Value: %h\n", PRED44_11_buffer[clk]);
        end
        if (PRED44_12_buffer[clk] != PRED44_12_buffer[!clk]) begin
          $fwrite(f, "Register (44,12) Value: %h\n", PRED44_12_buffer[clk]);
        end
        if (PRED44_13_buffer[clk] != PRED44_13_buffer[!clk]) begin
          $fwrite(f, "Register (44,13) Value: %h\n", PRED44_13_buffer[clk]);
        end
        if (PRED44_14_buffer[clk] != PRED44_14_buffer[!clk]) begin
          $fwrite(f, "Register (44,14) Value: %h\n", PRED44_14_buffer[clk]);
        end
        if (PRED44_15_buffer[clk] != PRED44_15_buffer[!clk]) begin
          $fwrite(f, "Register (44,15) Value: %h\n", PRED44_15_buffer[clk]);
        end
        if (PRED44_16_buffer[clk] != PRED44_16_buffer[!clk]) begin
          $fwrite(f, "Register (44,16) Value: %h\n", PRED44_16_buffer[clk]);
        end
        if (PRED44_17_buffer[clk] != PRED44_17_buffer[!clk]) begin
          $fwrite(f, "Register (44,17) Value: %h\n", PRED44_17_buffer[clk]);
        end
        if (PRED44_18_buffer[clk] != PRED44_18_buffer[!clk]) begin
          $fwrite(f, "Register (44,18) Value: %h\n", PRED44_18_buffer[clk]);
        end
        if (PRED44_19_buffer[clk] != PRED44_19_buffer[!clk]) begin
          $fwrite(f, "Register (44,19) Value: %h\n", PRED44_19_buffer[clk]);
        end
        if (PRED44_20_buffer[clk] != PRED44_20_buffer[!clk]) begin
          $fwrite(f, "Register (44,20) Value: %h\n", PRED44_20_buffer[clk]);
        end
        if (PRED44_21_buffer[clk] != PRED44_21_buffer[!clk]) begin
          $fwrite(f, "Register (44,21) Value: %h\n", PRED44_21_buffer[clk]);
        end
        if (PRED44_22_buffer[clk] != PRED44_22_buffer[!clk]) begin
          $fwrite(f, "Register (44,22) Value: %h\n", PRED44_22_buffer[clk]);
        end
        if (PRED44_23_buffer[clk] != PRED44_23_buffer[!clk]) begin
          $fwrite(f, "Register (44,23) Value: %h\n", PRED44_23_buffer[clk]);
        end
        if (PRED44_24_buffer[clk] != PRED44_24_buffer[!clk]) begin
          $fwrite(f, "Register (44,24) Value: %h\n", PRED44_24_buffer[clk]);
        end
        if (PRED44_25_buffer[clk] != PRED44_25_buffer[!clk]) begin
          $fwrite(f, "Register (44,25) Value: %h\n", PRED44_25_buffer[clk]);
        end
        if (PRED44_26_buffer[clk] != PRED44_26_buffer[!clk]) begin
          $fwrite(f, "Register (44,26) Value: %h\n", PRED44_26_buffer[clk]);
        end
        if (PRED44_27_buffer[clk] != PRED44_27_buffer[!clk]) begin
          $fwrite(f, "Register (44,27) Value: %h\n", PRED44_27_buffer[clk]);
        end
        if (PRED44_28_buffer[clk] != PRED44_28_buffer[!clk]) begin
          $fwrite(f, "Register (44,28) Value: %h\n", PRED44_28_buffer[clk]);
        end
        if (PRED44_29_buffer[clk] != PRED44_29_buffer[!clk]) begin
          $fwrite(f, "Register (44,29) Value: %h\n", PRED44_29_buffer[clk]);
        end
        if (PRED44_30_buffer[clk] != PRED44_30_buffer[!clk]) begin
          $fwrite(f, "Register (44,30) Value: %h\n", PRED44_30_buffer[clk]);
        end
        if (PRED44_31_buffer[clk] != PRED44_31_buffer[!clk]) begin
          $fwrite(f, "Register (44,31) Value: %h\n", PRED44_31_buffer[clk]);
        end
        if (PRED45_0_buffer[clk] != PRED45_0_buffer[!clk]) begin
          $fwrite(f, "Register (45,0) Value: %h\n", PRED45_0_buffer[clk]);
        end
        if (PRED45_1_buffer[clk] != PRED45_1_buffer[!clk]) begin
          $fwrite(f, "Register (45,1) Value: %h\n", PRED45_1_buffer[clk]);
        end
        if (PRED45_2_buffer[clk] != PRED45_2_buffer[!clk]) begin
          $fwrite(f, "Register (45,2) Value: %h\n", PRED45_2_buffer[clk]);
        end
        if (PRED45_3_buffer[clk] != PRED45_3_buffer[!clk]) begin
          $fwrite(f, "Register (45,3) Value: %h\n", PRED45_3_buffer[clk]);
        end
        if (PRED45_4_buffer[clk] != PRED45_4_buffer[!clk]) begin
          $fwrite(f, "Register (45,4) Value: %h\n", PRED45_4_buffer[clk]);
        end
        if (PRED45_5_buffer[clk] != PRED45_5_buffer[!clk]) begin
          $fwrite(f, "Register (45,5) Value: %h\n", PRED45_5_buffer[clk]);
        end
        if (PRED45_6_buffer[clk] != PRED45_6_buffer[!clk]) begin
          $fwrite(f, "Register (45,6) Value: %h\n", PRED45_6_buffer[clk]);
        end
        if (PRED45_7_buffer[clk] != PRED45_7_buffer[!clk]) begin
          $fwrite(f, "Register (45,7) Value: %h\n", PRED45_7_buffer[clk]);
        end
        if (PRED45_8_buffer[clk] != PRED45_8_buffer[!clk]) begin
          $fwrite(f, "Register (45,8) Value: %h\n", PRED45_8_buffer[clk]);
        end
        if (PRED45_9_buffer[clk] != PRED45_9_buffer[!clk]) begin
          $fwrite(f, "Register (45,9) Value: %h\n", PRED45_9_buffer[clk]);
        end
        if (PRED45_10_buffer[clk] != PRED45_10_buffer[!clk]) begin
          $fwrite(f, "Register (45,10) Value: %h\n", PRED45_10_buffer[clk]);
        end
        if (PRED45_11_buffer[clk] != PRED45_11_buffer[!clk]) begin
          $fwrite(f, "Register (45,11) Value: %h\n", PRED45_11_buffer[clk]);
        end
        if (PRED45_12_buffer[clk] != PRED45_12_buffer[!clk]) begin
          $fwrite(f, "Register (45,12) Value: %h\n", PRED45_12_buffer[clk]);
        end
        if (PRED45_13_buffer[clk] != PRED45_13_buffer[!clk]) begin
          $fwrite(f, "Register (45,13) Value: %h\n", PRED45_13_buffer[clk]);
        end
        if (PRED45_14_buffer[clk] != PRED45_14_buffer[!clk]) begin
          $fwrite(f, "Register (45,14) Value: %h\n", PRED45_14_buffer[clk]);
        end
        if (PRED45_15_buffer[clk] != PRED45_15_buffer[!clk]) begin
          $fwrite(f, "Register (45,15) Value: %h\n", PRED45_15_buffer[clk]);
        end
        if (PRED45_16_buffer[clk] != PRED45_16_buffer[!clk]) begin
          $fwrite(f, "Register (45,16) Value: %h\n", PRED45_16_buffer[clk]);
        end
        if (PRED45_17_buffer[clk] != PRED45_17_buffer[!clk]) begin
          $fwrite(f, "Register (45,17) Value: %h\n", PRED45_17_buffer[clk]);
        end
        if (PRED45_18_buffer[clk] != PRED45_18_buffer[!clk]) begin
          $fwrite(f, "Register (45,18) Value: %h\n", PRED45_18_buffer[clk]);
        end
        if (PRED45_19_buffer[clk] != PRED45_19_buffer[!clk]) begin
          $fwrite(f, "Register (45,19) Value: %h\n", PRED45_19_buffer[clk]);
        end
        if (PRED45_20_buffer[clk] != PRED45_20_buffer[!clk]) begin
          $fwrite(f, "Register (45,20) Value: %h\n", PRED45_20_buffer[clk]);
        end
        if (PRED45_21_buffer[clk] != PRED45_21_buffer[!clk]) begin
          $fwrite(f, "Register (45,21) Value: %h\n", PRED45_21_buffer[clk]);
        end
        if (PRED45_22_buffer[clk] != PRED45_22_buffer[!clk]) begin
          $fwrite(f, "Register (45,22) Value: %h\n", PRED45_22_buffer[clk]);
        end
        if (PRED45_23_buffer[clk] != PRED45_23_buffer[!clk]) begin
          $fwrite(f, "Register (45,23) Value: %h\n", PRED45_23_buffer[clk]);
        end
        if (PRED45_24_buffer[clk] != PRED45_24_buffer[!clk]) begin
          $fwrite(f, "Register (45,24) Value: %h\n", PRED45_24_buffer[clk]);
        end
        if (PRED45_25_buffer[clk] != PRED45_25_buffer[!clk]) begin
          $fwrite(f, "Register (45,25) Value: %h\n", PRED45_25_buffer[clk]);
        end
        if (PRED45_26_buffer[clk] != PRED45_26_buffer[!clk]) begin
          $fwrite(f, "Register (45,26) Value: %h\n", PRED45_26_buffer[clk]);
        end
        if (PRED45_27_buffer[clk] != PRED45_27_buffer[!clk]) begin
          $fwrite(f, "Register (45,27) Value: %h\n", PRED45_27_buffer[clk]);
        end
        if (PRED45_28_buffer[clk] != PRED45_28_buffer[!clk]) begin
          $fwrite(f, "Register (45,28) Value: %h\n", PRED45_28_buffer[clk]);
        end
        if (PRED45_29_buffer[clk] != PRED45_29_buffer[!clk]) begin
          $fwrite(f, "Register (45,29) Value: %h\n", PRED45_29_buffer[clk]);
        end
        if (PRED45_30_buffer[clk] != PRED45_30_buffer[!clk]) begin
          $fwrite(f, "Register (45,30) Value: %h\n", PRED45_30_buffer[clk]);
        end
        if (PRED45_31_buffer[clk] != PRED45_31_buffer[!clk]) begin
          $fwrite(f, "Register (45,31) Value: %h\n", PRED45_31_buffer[clk]);
        end
        if (PRED46_0_buffer[clk] != PRED46_0_buffer[!clk]) begin
          $fwrite(f, "Register (46,0) Value: %h\n", PRED46_0_buffer[clk]);
        end
        if (PRED46_1_buffer[clk] != PRED46_1_buffer[!clk]) begin
          $fwrite(f, "Register (46,1) Value: %h\n", PRED46_1_buffer[clk]);
        end
        if (PRED46_2_buffer[clk] != PRED46_2_buffer[!clk]) begin
          $fwrite(f, "Register (46,2) Value: %h\n", PRED46_2_buffer[clk]);
        end
        if (PRED46_3_buffer[clk] != PRED46_3_buffer[!clk]) begin
          $fwrite(f, "Register (46,3) Value: %h\n", PRED46_3_buffer[clk]);
        end
        if (PRED46_4_buffer[clk] != PRED46_4_buffer[!clk]) begin
          $fwrite(f, "Register (46,4) Value: %h\n", PRED46_4_buffer[clk]);
        end
        if (PRED46_5_buffer[clk] != PRED46_5_buffer[!clk]) begin
          $fwrite(f, "Register (46,5) Value: %h\n", PRED46_5_buffer[clk]);
        end
        if (PRED46_6_buffer[clk] != PRED46_6_buffer[!clk]) begin
          $fwrite(f, "Register (46,6) Value: %h\n", PRED46_6_buffer[clk]);
        end
        if (PRED46_7_buffer[clk] != PRED46_7_buffer[!clk]) begin
          $fwrite(f, "Register (46,7) Value: %h\n", PRED46_7_buffer[clk]);
        end
        if (PRED46_8_buffer[clk] != PRED46_8_buffer[!clk]) begin
          $fwrite(f, "Register (46,8) Value: %h\n", PRED46_8_buffer[clk]);
        end
        if (PRED46_9_buffer[clk] != PRED46_9_buffer[!clk]) begin
          $fwrite(f, "Register (46,9) Value: %h\n", PRED46_9_buffer[clk]);
        end
        if (PRED46_10_buffer[clk] != PRED46_10_buffer[!clk]) begin
          $fwrite(f, "Register (46,10) Value: %h\n", PRED46_10_buffer[clk]);
        end
        if (PRED46_11_buffer[clk] != PRED46_11_buffer[!clk]) begin
          $fwrite(f, "Register (46,11) Value: %h\n", PRED46_11_buffer[clk]);
        end
        if (PRED46_12_buffer[clk] != PRED46_12_buffer[!clk]) begin
          $fwrite(f, "Register (46,12) Value: %h\n", PRED46_12_buffer[clk]);
        end
        if (PRED46_13_buffer[clk] != PRED46_13_buffer[!clk]) begin
          $fwrite(f, "Register (46,13) Value: %h\n", PRED46_13_buffer[clk]);
        end
        if (PRED46_14_buffer[clk] != PRED46_14_buffer[!clk]) begin
          $fwrite(f, "Register (46,14) Value: %h\n", PRED46_14_buffer[clk]);
        end
        if (PRED46_15_buffer[clk] != PRED46_15_buffer[!clk]) begin
          $fwrite(f, "Register (46,15) Value: %h\n", PRED46_15_buffer[clk]);
        end
        if (PRED46_16_buffer[clk] != PRED46_16_buffer[!clk]) begin
          $fwrite(f, "Register (46,16) Value: %h\n", PRED46_16_buffer[clk]);
        end
        if (PRED46_17_buffer[clk] != PRED46_17_buffer[!clk]) begin
          $fwrite(f, "Register (46,17) Value: %h\n", PRED46_17_buffer[clk]);
        end
        if (PRED46_18_buffer[clk] != PRED46_18_buffer[!clk]) begin
          $fwrite(f, "Register (46,18) Value: %h\n", PRED46_18_buffer[clk]);
        end
        if (PRED46_19_buffer[clk] != PRED46_19_buffer[!clk]) begin
          $fwrite(f, "Register (46,19) Value: %h\n", PRED46_19_buffer[clk]);
        end
        if (PRED46_20_buffer[clk] != PRED46_20_buffer[!clk]) begin
          $fwrite(f, "Register (46,20) Value: %h\n", PRED46_20_buffer[clk]);
        end
        if (PRED46_21_buffer[clk] != PRED46_21_buffer[!clk]) begin
          $fwrite(f, "Register (46,21) Value: %h\n", PRED46_21_buffer[clk]);
        end
        if (PRED46_22_buffer[clk] != PRED46_22_buffer[!clk]) begin
          $fwrite(f, "Register (46,22) Value: %h\n", PRED46_22_buffer[clk]);
        end
        if (PRED46_23_buffer[clk] != PRED46_23_buffer[!clk]) begin
          $fwrite(f, "Register (46,23) Value: %h\n", PRED46_23_buffer[clk]);
        end
        if (PRED46_24_buffer[clk] != PRED46_24_buffer[!clk]) begin
          $fwrite(f, "Register (46,24) Value: %h\n", PRED46_24_buffer[clk]);
        end
        if (PRED46_25_buffer[clk] != PRED46_25_buffer[!clk]) begin
          $fwrite(f, "Register (46,25) Value: %h\n", PRED46_25_buffer[clk]);
        end
        if (PRED46_26_buffer[clk] != PRED46_26_buffer[!clk]) begin
          $fwrite(f, "Register (46,26) Value: %h\n", PRED46_26_buffer[clk]);
        end
        if (PRED46_27_buffer[clk] != PRED46_27_buffer[!clk]) begin
          $fwrite(f, "Register (46,27) Value: %h\n", PRED46_27_buffer[clk]);
        end
        if (PRED46_28_buffer[clk] != PRED46_28_buffer[!clk]) begin
          $fwrite(f, "Register (46,28) Value: %h\n", PRED46_28_buffer[clk]);
        end
        if (PRED46_29_buffer[clk] != PRED46_29_buffer[!clk]) begin
          $fwrite(f, "Register (46,29) Value: %h\n", PRED46_29_buffer[clk]);
        end
        if (PRED46_30_buffer[clk] != PRED46_30_buffer[!clk]) begin
          $fwrite(f, "Register (46,30) Value: %h\n", PRED46_30_buffer[clk]);
        end
        if (PRED46_31_buffer[clk] != PRED46_31_buffer[!clk]) begin
          $fwrite(f, "Register (46,31) Value: %h\n", PRED46_31_buffer[clk]);
        end
        if (PRED47_0_buffer[clk] != PRED47_0_buffer[!clk]) begin
          $fwrite(f, "Register (47,0) Value: %h\n", PRED47_0_buffer[clk]);
        end
        if (PRED47_1_buffer[clk] != PRED47_1_buffer[!clk]) begin
          $fwrite(f, "Register (47,1) Value: %h\n", PRED47_1_buffer[clk]);
        end
        if (PRED47_2_buffer[clk] != PRED47_2_buffer[!clk]) begin
          $fwrite(f, "Register (47,2) Value: %h\n", PRED47_2_buffer[clk]);
        end
        if (PRED47_3_buffer[clk] != PRED47_3_buffer[!clk]) begin
          $fwrite(f, "Register (47,3) Value: %h\n", PRED47_3_buffer[clk]);
        end
        if (PRED47_4_buffer[clk] != PRED47_4_buffer[!clk]) begin
          $fwrite(f, "Register (47,4) Value: %h\n", PRED47_4_buffer[clk]);
        end
        if (PRED47_5_buffer[clk] != PRED47_5_buffer[!clk]) begin
          $fwrite(f, "Register (47,5) Value: %h\n", PRED47_5_buffer[clk]);
        end
        if (PRED47_6_buffer[clk] != PRED47_6_buffer[!clk]) begin
          $fwrite(f, "Register (47,6) Value: %h\n", PRED47_6_buffer[clk]);
        end
        if (PRED47_7_buffer[clk] != PRED47_7_buffer[!clk]) begin
          $fwrite(f, "Register (47,7) Value: %h\n", PRED47_7_buffer[clk]);
        end
        if (PRED47_8_buffer[clk] != PRED47_8_buffer[!clk]) begin
          $fwrite(f, "Register (47,8) Value: %h\n", PRED47_8_buffer[clk]);
        end
        if (PRED47_9_buffer[clk] != PRED47_9_buffer[!clk]) begin
          $fwrite(f, "Register (47,9) Value: %h\n", PRED47_9_buffer[clk]);
        end
        if (PRED47_10_buffer[clk] != PRED47_10_buffer[!clk]) begin
          $fwrite(f, "Register (47,10) Value: %h\n", PRED47_10_buffer[clk]);
        end
        if (PRED47_11_buffer[clk] != PRED47_11_buffer[!clk]) begin
          $fwrite(f, "Register (47,11) Value: %h\n", PRED47_11_buffer[clk]);
        end
        if (PRED47_12_buffer[clk] != PRED47_12_buffer[!clk]) begin
          $fwrite(f, "Register (47,12) Value: %h\n", PRED47_12_buffer[clk]);
        end
        if (PRED47_13_buffer[clk] != PRED47_13_buffer[!clk]) begin
          $fwrite(f, "Register (47,13) Value: %h\n", PRED47_13_buffer[clk]);
        end
        if (PRED47_14_buffer[clk] != PRED47_14_buffer[!clk]) begin
          $fwrite(f, "Register (47,14) Value: %h\n", PRED47_14_buffer[clk]);
        end
        if (PRED47_15_buffer[clk] != PRED47_15_buffer[!clk]) begin
          $fwrite(f, "Register (47,15) Value: %h\n", PRED47_15_buffer[clk]);
        end
        if (PRED47_16_buffer[clk] != PRED47_16_buffer[!clk]) begin
          $fwrite(f, "Register (47,16) Value: %h\n", PRED47_16_buffer[clk]);
        end
        if (PRED47_17_buffer[clk] != PRED47_17_buffer[!clk]) begin
          $fwrite(f, "Register (47,17) Value: %h\n", PRED47_17_buffer[clk]);
        end
        if (PRED47_18_buffer[clk] != PRED47_18_buffer[!clk]) begin
          $fwrite(f, "Register (47,18) Value: %h\n", PRED47_18_buffer[clk]);
        end
        if (PRED47_19_buffer[clk] != PRED47_19_buffer[!clk]) begin
          $fwrite(f, "Register (47,19) Value: %h\n", PRED47_19_buffer[clk]);
        end
        if (PRED47_20_buffer[clk] != PRED47_20_buffer[!clk]) begin
          $fwrite(f, "Register (47,20) Value: %h\n", PRED47_20_buffer[clk]);
        end
        if (PRED47_21_buffer[clk] != PRED47_21_buffer[!clk]) begin
          $fwrite(f, "Register (47,21) Value: %h\n", PRED47_21_buffer[clk]);
        end
        if (PRED47_22_buffer[clk] != PRED47_22_buffer[!clk]) begin
          $fwrite(f, "Register (47,22) Value: %h\n", PRED47_22_buffer[clk]);
        end
        if (PRED47_23_buffer[clk] != PRED47_23_buffer[!clk]) begin
          $fwrite(f, "Register (47,23) Value: %h\n", PRED47_23_buffer[clk]);
        end
        if (PRED47_24_buffer[clk] != PRED47_24_buffer[!clk]) begin
          $fwrite(f, "Register (47,24) Value: %h\n", PRED47_24_buffer[clk]);
        end
        if (PRED47_25_buffer[clk] != PRED47_25_buffer[!clk]) begin
          $fwrite(f, "Register (47,25) Value: %h\n", PRED47_25_buffer[clk]);
        end
        if (PRED47_26_buffer[clk] != PRED47_26_buffer[!clk]) begin
          $fwrite(f, "Register (47,26) Value: %h\n", PRED47_26_buffer[clk]);
        end
        if (PRED47_27_buffer[clk] != PRED47_27_buffer[!clk]) begin
          $fwrite(f, "Register (47,27) Value: %h\n", PRED47_27_buffer[clk]);
        end
        if (PRED47_28_buffer[clk] != PRED47_28_buffer[!clk]) begin
          $fwrite(f, "Register (47,28) Value: %h\n", PRED47_28_buffer[clk]);
        end
        if (PRED47_29_buffer[clk] != PRED47_29_buffer[!clk]) begin
          $fwrite(f, "Register (47,29) Value: %h\n", PRED47_29_buffer[clk]);
        end
        if (PRED47_30_buffer[clk] != PRED47_30_buffer[!clk]) begin
          $fwrite(f, "Register (47,30) Value: %h\n", PRED47_30_buffer[clk]);
        end
        if (PRED47_31_buffer[clk] != PRED47_31_buffer[!clk]) begin
          $fwrite(f, "Register (47,31) Value: %h\n", PRED47_31_buffer[clk]);
        end
        if (PRED48_0_buffer[clk] != PRED48_0_buffer[!clk]) begin
          $fwrite(f, "Register (48,0) Value: %h\n", PRED48_0_buffer[clk]);
        end
        if (PRED48_1_buffer[clk] != PRED48_1_buffer[!clk]) begin
          $fwrite(f, "Register (48,1) Value: %h\n", PRED48_1_buffer[clk]);
        end
        if (PRED48_2_buffer[clk] != PRED48_2_buffer[!clk]) begin
          $fwrite(f, "Register (48,2) Value: %h\n", PRED48_2_buffer[clk]);
        end
        if (PRED48_3_buffer[clk] != PRED48_3_buffer[!clk]) begin
          $fwrite(f, "Register (48,3) Value: %h\n", PRED48_3_buffer[clk]);
        end
        if (PRED48_4_buffer[clk] != PRED48_4_buffer[!clk]) begin
          $fwrite(f, "Register (48,4) Value: %h\n", PRED48_4_buffer[clk]);
        end
        if (PRED48_5_buffer[clk] != PRED48_5_buffer[!clk]) begin
          $fwrite(f, "Register (48,5) Value: %h\n", PRED48_5_buffer[clk]);
        end
        if (PRED48_6_buffer[clk] != PRED48_6_buffer[!clk]) begin
          $fwrite(f, "Register (48,6) Value: %h\n", PRED48_6_buffer[clk]);
        end
        if (PRED48_7_buffer[clk] != PRED48_7_buffer[!clk]) begin
          $fwrite(f, "Register (48,7) Value: %h\n", PRED48_7_buffer[clk]);
        end
        if (PRED48_8_buffer[clk] != PRED48_8_buffer[!clk]) begin
          $fwrite(f, "Register (48,8) Value: %h\n", PRED48_8_buffer[clk]);
        end
        if (PRED48_9_buffer[clk] != PRED48_9_buffer[!clk]) begin
          $fwrite(f, "Register (48,9) Value: %h\n", PRED48_9_buffer[clk]);
        end
        if (PRED48_10_buffer[clk] != PRED48_10_buffer[!clk]) begin
          $fwrite(f, "Register (48,10) Value: %h\n", PRED48_10_buffer[clk]);
        end
        if (PRED48_11_buffer[clk] != PRED48_11_buffer[!clk]) begin
          $fwrite(f, "Register (48,11) Value: %h\n", PRED48_11_buffer[clk]);
        end
        if (PRED48_12_buffer[clk] != PRED48_12_buffer[!clk]) begin
          $fwrite(f, "Register (48,12) Value: %h\n", PRED48_12_buffer[clk]);
        end
        if (PRED48_13_buffer[clk] != PRED48_13_buffer[!clk]) begin
          $fwrite(f, "Register (48,13) Value: %h\n", PRED48_13_buffer[clk]);
        end
        if (PRED48_14_buffer[clk] != PRED48_14_buffer[!clk]) begin
          $fwrite(f, "Register (48,14) Value: %h\n", PRED48_14_buffer[clk]);
        end
        if (PRED48_15_buffer[clk] != PRED48_15_buffer[!clk]) begin
          $fwrite(f, "Register (48,15) Value: %h\n", PRED48_15_buffer[clk]);
        end
        if (PRED48_16_buffer[clk] != PRED48_16_buffer[!clk]) begin
          $fwrite(f, "Register (48,16) Value: %h\n", PRED48_16_buffer[clk]);
        end
        if (PRED48_17_buffer[clk] != PRED48_17_buffer[!clk]) begin
          $fwrite(f, "Register (48,17) Value: %h\n", PRED48_17_buffer[clk]);
        end
        if (PRED48_18_buffer[clk] != PRED48_18_buffer[!clk]) begin
          $fwrite(f, "Register (48,18) Value: %h\n", PRED48_18_buffer[clk]);
        end
        if (PRED48_19_buffer[clk] != PRED48_19_buffer[!clk]) begin
          $fwrite(f, "Register (48,19) Value: %h\n", PRED48_19_buffer[clk]);
        end
        if (PRED48_20_buffer[clk] != PRED48_20_buffer[!clk]) begin
          $fwrite(f, "Register (48,20) Value: %h\n", PRED48_20_buffer[clk]);
        end
        if (PRED48_21_buffer[clk] != PRED48_21_buffer[!clk]) begin
          $fwrite(f, "Register (48,21) Value: %h\n", PRED48_21_buffer[clk]);
        end
        if (PRED48_22_buffer[clk] != PRED48_22_buffer[!clk]) begin
          $fwrite(f, "Register (48,22) Value: %h\n", PRED48_22_buffer[clk]);
        end
        if (PRED48_23_buffer[clk] != PRED48_23_buffer[!clk]) begin
          $fwrite(f, "Register (48,23) Value: %h\n", PRED48_23_buffer[clk]);
        end
        if (PRED48_24_buffer[clk] != PRED48_24_buffer[!clk]) begin
          $fwrite(f, "Register (48,24) Value: %h\n", PRED48_24_buffer[clk]);
        end
        if (PRED48_25_buffer[clk] != PRED48_25_buffer[!clk]) begin
          $fwrite(f, "Register (48,25) Value: %h\n", PRED48_25_buffer[clk]);
        end
        if (PRED48_26_buffer[clk] != PRED48_26_buffer[!clk]) begin
          $fwrite(f, "Register (48,26) Value: %h\n", PRED48_26_buffer[clk]);
        end
        if (PRED48_27_buffer[clk] != PRED48_27_buffer[!clk]) begin
          $fwrite(f, "Register (48,27) Value: %h\n", PRED48_27_buffer[clk]);
        end
        if (PRED48_28_buffer[clk] != PRED48_28_buffer[!clk]) begin
          $fwrite(f, "Register (48,28) Value: %h\n", PRED48_28_buffer[clk]);
        end
        if (PRED48_29_buffer[clk] != PRED48_29_buffer[!clk]) begin
          $fwrite(f, "Register (48,29) Value: %h\n", PRED48_29_buffer[clk]);
        end
        if (PRED48_30_buffer[clk] != PRED48_30_buffer[!clk]) begin
          $fwrite(f, "Register (48,30) Value: %h\n", PRED48_30_buffer[clk]);
        end
        if (PRED48_31_buffer[clk] != PRED48_31_buffer[!clk]) begin
          $fwrite(f, "Register (48,31) Value: %h\n", PRED48_31_buffer[clk]);
        end
        if (PRED49_0_buffer[clk] != PRED49_0_buffer[!clk]) begin
          $fwrite(f, "Register (49,0) Value: %h\n", PRED49_0_buffer[clk]);
        end
        if (PRED49_1_buffer[clk] != PRED49_1_buffer[!clk]) begin
          $fwrite(f, "Register (49,1) Value: %h\n", PRED49_1_buffer[clk]);
        end
        if (PRED49_2_buffer[clk] != PRED49_2_buffer[!clk]) begin
          $fwrite(f, "Register (49,2) Value: %h\n", PRED49_2_buffer[clk]);
        end
        if (PRED49_3_buffer[clk] != PRED49_3_buffer[!clk]) begin
          $fwrite(f, "Register (49,3) Value: %h\n", PRED49_3_buffer[clk]);
        end
        if (PRED49_4_buffer[clk] != PRED49_4_buffer[!clk]) begin
          $fwrite(f, "Register (49,4) Value: %h\n", PRED49_4_buffer[clk]);
        end
        if (PRED49_5_buffer[clk] != PRED49_5_buffer[!clk]) begin
          $fwrite(f, "Register (49,5) Value: %h\n", PRED49_5_buffer[clk]);
        end
        if (PRED49_6_buffer[clk] != PRED49_6_buffer[!clk]) begin
          $fwrite(f, "Register (49,6) Value: %h\n", PRED49_6_buffer[clk]);
        end
        if (PRED49_7_buffer[clk] != PRED49_7_buffer[!clk]) begin
          $fwrite(f, "Register (49,7) Value: %h\n", PRED49_7_buffer[clk]);
        end
        if (PRED49_8_buffer[clk] != PRED49_8_buffer[!clk]) begin
          $fwrite(f, "Register (49,8) Value: %h\n", PRED49_8_buffer[clk]);
        end
        if (PRED49_9_buffer[clk] != PRED49_9_buffer[!clk]) begin
          $fwrite(f, "Register (49,9) Value: %h\n", PRED49_9_buffer[clk]);
        end
        if (PRED49_10_buffer[clk] != PRED49_10_buffer[!clk]) begin
          $fwrite(f, "Register (49,10) Value: %h\n", PRED49_10_buffer[clk]);
        end
        if (PRED49_11_buffer[clk] != PRED49_11_buffer[!clk]) begin
          $fwrite(f, "Register (49,11) Value: %h\n", PRED49_11_buffer[clk]);
        end
        if (PRED49_12_buffer[clk] != PRED49_12_buffer[!clk]) begin
          $fwrite(f, "Register (49,12) Value: %h\n", PRED49_12_buffer[clk]);
        end
        if (PRED49_13_buffer[clk] != PRED49_13_buffer[!clk]) begin
          $fwrite(f, "Register (49,13) Value: %h\n", PRED49_13_buffer[clk]);
        end
        if (PRED49_14_buffer[clk] != PRED49_14_buffer[!clk]) begin
          $fwrite(f, "Register (49,14) Value: %h\n", PRED49_14_buffer[clk]);
        end
        if (PRED49_15_buffer[clk] != PRED49_15_buffer[!clk]) begin
          $fwrite(f, "Register (49,15) Value: %h\n", PRED49_15_buffer[clk]);
        end
        if (PRED49_16_buffer[clk] != PRED49_16_buffer[!clk]) begin
          $fwrite(f, "Register (49,16) Value: %h\n", PRED49_16_buffer[clk]);
        end
        if (PRED49_17_buffer[clk] != PRED49_17_buffer[!clk]) begin
          $fwrite(f, "Register (49,17) Value: %h\n", PRED49_17_buffer[clk]);
        end
        if (PRED49_18_buffer[clk] != PRED49_18_buffer[!clk]) begin
          $fwrite(f, "Register (49,18) Value: %h\n", PRED49_18_buffer[clk]);
        end
        if (PRED49_19_buffer[clk] != PRED49_19_buffer[!clk]) begin
          $fwrite(f, "Register (49,19) Value: %h\n", PRED49_19_buffer[clk]);
        end
        if (PRED49_20_buffer[clk] != PRED49_20_buffer[!clk]) begin
          $fwrite(f, "Register (49,20) Value: %h\n", PRED49_20_buffer[clk]);
        end
        if (PRED49_21_buffer[clk] != PRED49_21_buffer[!clk]) begin
          $fwrite(f, "Register (49,21) Value: %h\n", PRED49_21_buffer[clk]);
        end
        if (PRED49_22_buffer[clk] != PRED49_22_buffer[!clk]) begin
          $fwrite(f, "Register (49,22) Value: %h\n", PRED49_22_buffer[clk]);
        end
        if (PRED49_23_buffer[clk] != PRED49_23_buffer[!clk]) begin
          $fwrite(f, "Register (49,23) Value: %h\n", PRED49_23_buffer[clk]);
        end
        if (PRED49_24_buffer[clk] != PRED49_24_buffer[!clk]) begin
          $fwrite(f, "Register (49,24) Value: %h\n", PRED49_24_buffer[clk]);
        end
        if (PRED49_25_buffer[clk] != PRED49_25_buffer[!clk]) begin
          $fwrite(f, "Register (49,25) Value: %h\n", PRED49_25_buffer[clk]);
        end
        if (PRED49_26_buffer[clk] != PRED49_26_buffer[!clk]) begin
          $fwrite(f, "Register (49,26) Value: %h\n", PRED49_26_buffer[clk]);
        end
        if (PRED49_27_buffer[clk] != PRED49_27_buffer[!clk]) begin
          $fwrite(f, "Register (49,27) Value: %h\n", PRED49_27_buffer[clk]);
        end
        if (PRED49_28_buffer[clk] != PRED49_28_buffer[!clk]) begin
          $fwrite(f, "Register (49,28) Value: %h\n", PRED49_28_buffer[clk]);
        end
        if (PRED49_29_buffer[clk] != PRED49_29_buffer[!clk]) begin
          $fwrite(f, "Register (49,29) Value: %h\n", PRED49_29_buffer[clk]);
        end
        if (PRED49_30_buffer[clk] != PRED49_30_buffer[!clk]) begin
          $fwrite(f, "Register (49,30) Value: %h\n", PRED49_30_buffer[clk]);
        end
        if (PRED49_31_buffer[clk] != PRED49_31_buffer[!clk]) begin
          $fwrite(f, "Register (49,31) Value: %h\n", PRED49_31_buffer[clk]);
        end
        if (PRED50_0_buffer[clk] != PRED50_0_buffer[!clk]) begin
          $fwrite(f, "Register (50,0) Value: %h\n", PRED50_0_buffer[clk]);
        end
        if (PRED50_1_buffer[clk] != PRED50_1_buffer[!clk]) begin
          $fwrite(f, "Register (50,1) Value: %h\n", PRED50_1_buffer[clk]);
        end
        if (PRED50_2_buffer[clk] != PRED50_2_buffer[!clk]) begin
          $fwrite(f, "Register (50,2) Value: %h\n", PRED50_2_buffer[clk]);
        end
        if (PRED50_3_buffer[clk] != PRED50_3_buffer[!clk]) begin
          $fwrite(f, "Register (50,3) Value: %h\n", PRED50_3_buffer[clk]);
        end
        if (PRED50_4_buffer[clk] != PRED50_4_buffer[!clk]) begin
          $fwrite(f, "Register (50,4) Value: %h\n", PRED50_4_buffer[clk]);
        end
        if (PRED50_5_buffer[clk] != PRED50_5_buffer[!clk]) begin
          $fwrite(f, "Register (50,5) Value: %h\n", PRED50_5_buffer[clk]);
        end
        if (PRED50_6_buffer[clk] != PRED50_6_buffer[!clk]) begin
          $fwrite(f, "Register (50,6) Value: %h\n", PRED50_6_buffer[clk]);
        end
        if (PRED50_7_buffer[clk] != PRED50_7_buffer[!clk]) begin
          $fwrite(f, "Register (50,7) Value: %h\n", PRED50_7_buffer[clk]);
        end
        if (PRED50_8_buffer[clk] != PRED50_8_buffer[!clk]) begin
          $fwrite(f, "Register (50,8) Value: %h\n", PRED50_8_buffer[clk]);
        end
        if (PRED50_9_buffer[clk] != PRED50_9_buffer[!clk]) begin
          $fwrite(f, "Register (50,9) Value: %h\n", PRED50_9_buffer[clk]);
        end
        if (PRED50_10_buffer[clk] != PRED50_10_buffer[!clk]) begin
          $fwrite(f, "Register (50,10) Value: %h\n", PRED50_10_buffer[clk]);
        end
        if (PRED50_11_buffer[clk] != PRED50_11_buffer[!clk]) begin
          $fwrite(f, "Register (50,11) Value: %h\n", PRED50_11_buffer[clk]);
        end
        if (PRED50_12_buffer[clk] != PRED50_12_buffer[!clk]) begin
          $fwrite(f, "Register (50,12) Value: %h\n", PRED50_12_buffer[clk]);
        end
        if (PRED50_13_buffer[clk] != PRED50_13_buffer[!clk]) begin
          $fwrite(f, "Register (50,13) Value: %h\n", PRED50_13_buffer[clk]);
        end
        if (PRED50_14_buffer[clk] != PRED50_14_buffer[!clk]) begin
          $fwrite(f, "Register (50,14) Value: %h\n", PRED50_14_buffer[clk]);
        end
        if (PRED50_15_buffer[clk] != PRED50_15_buffer[!clk]) begin
          $fwrite(f, "Register (50,15) Value: %h\n", PRED50_15_buffer[clk]);
        end
        if (PRED50_16_buffer[clk] != PRED50_16_buffer[!clk]) begin
          $fwrite(f, "Register (50,16) Value: %h\n", PRED50_16_buffer[clk]);
        end
        if (PRED50_17_buffer[clk] != PRED50_17_buffer[!clk]) begin
          $fwrite(f, "Register (50,17) Value: %h\n", PRED50_17_buffer[clk]);
        end
        if (PRED50_18_buffer[clk] != PRED50_18_buffer[!clk]) begin
          $fwrite(f, "Register (50,18) Value: %h\n", PRED50_18_buffer[clk]);
        end
        if (PRED50_19_buffer[clk] != PRED50_19_buffer[!clk]) begin
          $fwrite(f, "Register (50,19) Value: %h\n", PRED50_19_buffer[clk]);
        end
        if (PRED50_20_buffer[clk] != PRED50_20_buffer[!clk]) begin
          $fwrite(f, "Register (50,20) Value: %h\n", PRED50_20_buffer[clk]);
        end
        if (PRED50_21_buffer[clk] != PRED50_21_buffer[!clk]) begin
          $fwrite(f, "Register (50,21) Value: %h\n", PRED50_21_buffer[clk]);
        end
        if (PRED50_22_buffer[clk] != PRED50_22_buffer[!clk]) begin
          $fwrite(f, "Register (50,22) Value: %h\n", PRED50_22_buffer[clk]);
        end
        if (PRED50_23_buffer[clk] != PRED50_23_buffer[!clk]) begin
          $fwrite(f, "Register (50,23) Value: %h\n", PRED50_23_buffer[clk]);
        end
        if (PRED50_24_buffer[clk] != PRED50_24_buffer[!clk]) begin
          $fwrite(f, "Register (50,24) Value: %h\n", PRED50_24_buffer[clk]);
        end
        if (PRED50_25_buffer[clk] != PRED50_25_buffer[!clk]) begin
          $fwrite(f, "Register (50,25) Value: %h\n", PRED50_25_buffer[clk]);
        end
        if (PRED50_26_buffer[clk] != PRED50_26_buffer[!clk]) begin
          $fwrite(f, "Register (50,26) Value: %h\n", PRED50_26_buffer[clk]);
        end
        if (PRED50_27_buffer[clk] != PRED50_27_buffer[!clk]) begin
          $fwrite(f, "Register (50,27) Value: %h\n", PRED50_27_buffer[clk]);
        end
        if (PRED50_28_buffer[clk] != PRED50_28_buffer[!clk]) begin
          $fwrite(f, "Register (50,28) Value: %h\n", PRED50_28_buffer[clk]);
        end
        if (PRED50_29_buffer[clk] != PRED50_29_buffer[!clk]) begin
          $fwrite(f, "Register (50,29) Value: %h\n", PRED50_29_buffer[clk]);
        end
        if (PRED50_30_buffer[clk] != PRED50_30_buffer[!clk]) begin
          $fwrite(f, "Register (50,30) Value: %h\n", PRED50_30_buffer[clk]);
        end
        if (PRED50_31_buffer[clk] != PRED50_31_buffer[!clk]) begin
          $fwrite(f, "Register (50,31) Value: %h\n", PRED50_31_buffer[clk]);
        end
        if (PRED51_0_buffer[clk] != PRED51_0_buffer[!clk]) begin
          $fwrite(f, "Register (51,0) Value: %h\n", PRED51_0_buffer[clk]);
        end
        if (PRED51_1_buffer[clk] != PRED51_1_buffer[!clk]) begin
          $fwrite(f, "Register (51,1) Value: %h\n", PRED51_1_buffer[clk]);
        end
        if (PRED51_2_buffer[clk] != PRED51_2_buffer[!clk]) begin
          $fwrite(f, "Register (51,2) Value: %h\n", PRED51_2_buffer[clk]);
        end
        if (PRED51_3_buffer[clk] != PRED51_3_buffer[!clk]) begin
          $fwrite(f, "Register (51,3) Value: %h\n", PRED51_3_buffer[clk]);
        end
        if (PRED51_4_buffer[clk] != PRED51_4_buffer[!clk]) begin
          $fwrite(f, "Register (51,4) Value: %h\n", PRED51_4_buffer[clk]);
        end
        if (PRED51_5_buffer[clk] != PRED51_5_buffer[!clk]) begin
          $fwrite(f, "Register (51,5) Value: %h\n", PRED51_5_buffer[clk]);
        end
        if (PRED51_6_buffer[clk] != PRED51_6_buffer[!clk]) begin
          $fwrite(f, "Register (51,6) Value: %h\n", PRED51_6_buffer[clk]);
        end
        if (PRED51_7_buffer[clk] != PRED51_7_buffer[!clk]) begin
          $fwrite(f, "Register (51,7) Value: %h\n", PRED51_7_buffer[clk]);
        end
        if (PRED51_8_buffer[clk] != PRED51_8_buffer[!clk]) begin
          $fwrite(f, "Register (51,8) Value: %h\n", PRED51_8_buffer[clk]);
        end
        if (PRED51_9_buffer[clk] != PRED51_9_buffer[!clk]) begin
          $fwrite(f, "Register (51,9) Value: %h\n", PRED51_9_buffer[clk]);
        end
        if (PRED51_10_buffer[clk] != PRED51_10_buffer[!clk]) begin
          $fwrite(f, "Register (51,10) Value: %h\n", PRED51_10_buffer[clk]);
        end
        if (PRED51_11_buffer[clk] != PRED51_11_buffer[!clk]) begin
          $fwrite(f, "Register (51,11) Value: %h\n", PRED51_11_buffer[clk]);
        end
        if (PRED51_12_buffer[clk] != PRED51_12_buffer[!clk]) begin
          $fwrite(f, "Register (51,12) Value: %h\n", PRED51_12_buffer[clk]);
        end
        if (PRED51_13_buffer[clk] != PRED51_13_buffer[!clk]) begin
          $fwrite(f, "Register (51,13) Value: %h\n", PRED51_13_buffer[clk]);
        end
        if (PRED51_14_buffer[clk] != PRED51_14_buffer[!clk]) begin
          $fwrite(f, "Register (51,14) Value: %h\n", PRED51_14_buffer[clk]);
        end
        if (PRED51_15_buffer[clk] != PRED51_15_buffer[!clk]) begin
          $fwrite(f, "Register (51,15) Value: %h\n", PRED51_15_buffer[clk]);
        end
        if (PRED51_16_buffer[clk] != PRED51_16_buffer[!clk]) begin
          $fwrite(f, "Register (51,16) Value: %h\n", PRED51_16_buffer[clk]);
        end
        if (PRED51_17_buffer[clk] != PRED51_17_buffer[!clk]) begin
          $fwrite(f, "Register (51,17) Value: %h\n", PRED51_17_buffer[clk]);
        end
        if (PRED51_18_buffer[clk] != PRED51_18_buffer[!clk]) begin
          $fwrite(f, "Register (51,18) Value: %h\n", PRED51_18_buffer[clk]);
        end
        if (PRED51_19_buffer[clk] != PRED51_19_buffer[!clk]) begin
          $fwrite(f, "Register (51,19) Value: %h\n", PRED51_19_buffer[clk]);
        end
        if (PRED51_20_buffer[clk] != PRED51_20_buffer[!clk]) begin
          $fwrite(f, "Register (51,20) Value: %h\n", PRED51_20_buffer[clk]);
        end
        if (PRED51_21_buffer[clk] != PRED51_21_buffer[!clk]) begin
          $fwrite(f, "Register (51,21) Value: %h\n", PRED51_21_buffer[clk]);
        end
        if (PRED51_22_buffer[clk] != PRED51_22_buffer[!clk]) begin
          $fwrite(f, "Register (51,22) Value: %h\n", PRED51_22_buffer[clk]);
        end
        if (PRED51_23_buffer[clk] != PRED51_23_buffer[!clk]) begin
          $fwrite(f, "Register (51,23) Value: %h\n", PRED51_23_buffer[clk]);
        end
        if (PRED51_24_buffer[clk] != PRED51_24_buffer[!clk]) begin
          $fwrite(f, "Register (51,24) Value: %h\n", PRED51_24_buffer[clk]);
        end
        if (PRED51_25_buffer[clk] != PRED51_25_buffer[!clk]) begin
          $fwrite(f, "Register (51,25) Value: %h\n", PRED51_25_buffer[clk]);
        end
        if (PRED51_26_buffer[clk] != PRED51_26_buffer[!clk]) begin
          $fwrite(f, "Register (51,26) Value: %h\n", PRED51_26_buffer[clk]);
        end
        if (PRED51_27_buffer[clk] != PRED51_27_buffer[!clk]) begin
          $fwrite(f, "Register (51,27) Value: %h\n", PRED51_27_buffer[clk]);
        end
        if (PRED51_28_buffer[clk] != PRED51_28_buffer[!clk]) begin
          $fwrite(f, "Register (51,28) Value: %h\n", PRED51_28_buffer[clk]);
        end
        if (PRED51_29_buffer[clk] != PRED51_29_buffer[!clk]) begin
          $fwrite(f, "Register (51,29) Value: %h\n", PRED51_29_buffer[clk]);
        end
        if (PRED51_30_buffer[clk] != PRED51_30_buffer[!clk]) begin
          $fwrite(f, "Register (51,30) Value: %h\n", PRED51_30_buffer[clk]);
        end
        if (PRED51_31_buffer[clk] != PRED51_31_buffer[!clk]) begin
          $fwrite(f, "Register (51,31) Value: %h\n", PRED51_31_buffer[clk]);
        end
        if (PRED52_0_buffer[clk] != PRED52_0_buffer[!clk]) begin
          $fwrite(f, "Register (52,0) Value: %h\n", PRED52_0_buffer[clk]);
        end
        if (PRED52_1_buffer[clk] != PRED52_1_buffer[!clk]) begin
          $fwrite(f, "Register (52,1) Value: %h\n", PRED52_1_buffer[clk]);
        end
        if (PRED52_2_buffer[clk] != PRED52_2_buffer[!clk]) begin
          $fwrite(f, "Register (52,2) Value: %h\n", PRED52_2_buffer[clk]);
        end
        if (PRED52_3_buffer[clk] != PRED52_3_buffer[!clk]) begin
          $fwrite(f, "Register (52,3) Value: %h\n", PRED52_3_buffer[clk]);
        end
        if (PRED52_4_buffer[clk] != PRED52_4_buffer[!clk]) begin
          $fwrite(f, "Register (52,4) Value: %h\n", PRED52_4_buffer[clk]);
        end
        if (PRED52_5_buffer[clk] != PRED52_5_buffer[!clk]) begin
          $fwrite(f, "Register (52,5) Value: %h\n", PRED52_5_buffer[clk]);
        end
        if (PRED52_6_buffer[clk] != PRED52_6_buffer[!clk]) begin
          $fwrite(f, "Register (52,6) Value: %h\n", PRED52_6_buffer[clk]);
        end
        if (PRED52_7_buffer[clk] != PRED52_7_buffer[!clk]) begin
          $fwrite(f, "Register (52,7) Value: %h\n", PRED52_7_buffer[clk]);
        end
        if (PRED52_8_buffer[clk] != PRED52_8_buffer[!clk]) begin
          $fwrite(f, "Register (52,8) Value: %h\n", PRED52_8_buffer[clk]);
        end
        if (PRED52_9_buffer[clk] != PRED52_9_buffer[!clk]) begin
          $fwrite(f, "Register (52,9) Value: %h\n", PRED52_9_buffer[clk]);
        end
        if (PRED52_10_buffer[clk] != PRED52_10_buffer[!clk]) begin
          $fwrite(f, "Register (52,10) Value: %h\n", PRED52_10_buffer[clk]);
        end
        if (PRED52_11_buffer[clk] != PRED52_11_buffer[!clk]) begin
          $fwrite(f, "Register (52,11) Value: %h\n", PRED52_11_buffer[clk]);
        end
        if (PRED52_12_buffer[clk] != PRED52_12_buffer[!clk]) begin
          $fwrite(f, "Register (52,12) Value: %h\n", PRED52_12_buffer[clk]);
        end
        if (PRED52_13_buffer[clk] != PRED52_13_buffer[!clk]) begin
          $fwrite(f, "Register (52,13) Value: %h\n", PRED52_13_buffer[clk]);
        end
        if (PRED52_14_buffer[clk] != PRED52_14_buffer[!clk]) begin
          $fwrite(f, "Register (52,14) Value: %h\n", PRED52_14_buffer[clk]);
        end
        if (PRED52_15_buffer[clk] != PRED52_15_buffer[!clk]) begin
          $fwrite(f, "Register (52,15) Value: %h\n", PRED52_15_buffer[clk]);
        end
        if (PRED52_16_buffer[clk] != PRED52_16_buffer[!clk]) begin
          $fwrite(f, "Register (52,16) Value: %h\n", PRED52_16_buffer[clk]);
        end
        if (PRED52_17_buffer[clk] != PRED52_17_buffer[!clk]) begin
          $fwrite(f, "Register (52,17) Value: %h\n", PRED52_17_buffer[clk]);
        end
        if (PRED52_18_buffer[clk] != PRED52_18_buffer[!clk]) begin
          $fwrite(f, "Register (52,18) Value: %h\n", PRED52_18_buffer[clk]);
        end
        if (PRED52_19_buffer[clk] != PRED52_19_buffer[!clk]) begin
          $fwrite(f, "Register (52,19) Value: %h\n", PRED52_19_buffer[clk]);
        end
        if (PRED52_20_buffer[clk] != PRED52_20_buffer[!clk]) begin
          $fwrite(f, "Register (52,20) Value: %h\n", PRED52_20_buffer[clk]);
        end
        if (PRED52_21_buffer[clk] != PRED52_21_buffer[!clk]) begin
          $fwrite(f, "Register (52,21) Value: %h\n", PRED52_21_buffer[clk]);
        end
        if (PRED52_22_buffer[clk] != PRED52_22_buffer[!clk]) begin
          $fwrite(f, "Register (52,22) Value: %h\n", PRED52_22_buffer[clk]);
        end
        if (PRED52_23_buffer[clk] != PRED52_23_buffer[!clk]) begin
          $fwrite(f, "Register (52,23) Value: %h\n", PRED52_23_buffer[clk]);
        end
        if (PRED52_24_buffer[clk] != PRED52_24_buffer[!clk]) begin
          $fwrite(f, "Register (52,24) Value: %h\n", PRED52_24_buffer[clk]);
        end
        if (PRED52_25_buffer[clk] != PRED52_25_buffer[!clk]) begin
          $fwrite(f, "Register (52,25) Value: %h\n", PRED52_25_buffer[clk]);
        end
        if (PRED52_26_buffer[clk] != PRED52_26_buffer[!clk]) begin
          $fwrite(f, "Register (52,26) Value: %h\n", PRED52_26_buffer[clk]);
        end
        if (PRED52_27_buffer[clk] != PRED52_27_buffer[!clk]) begin
          $fwrite(f, "Register (52,27) Value: %h\n", PRED52_27_buffer[clk]);
        end
        if (PRED52_28_buffer[clk] != PRED52_28_buffer[!clk]) begin
          $fwrite(f, "Register (52,28) Value: %h\n", PRED52_28_buffer[clk]);
        end
        if (PRED52_29_buffer[clk] != PRED52_29_buffer[!clk]) begin
          $fwrite(f, "Register (52,29) Value: %h\n", PRED52_29_buffer[clk]);
        end
        if (PRED52_30_buffer[clk] != PRED52_30_buffer[!clk]) begin
          $fwrite(f, "Register (52,30) Value: %h\n", PRED52_30_buffer[clk]);
        end
        if (PRED52_31_buffer[clk] != PRED52_31_buffer[!clk]) begin
          $fwrite(f, "Register (52,31) Value: %h\n", PRED52_31_buffer[clk]);
        end
        if (PRED53_0_buffer[clk] != PRED53_0_buffer[!clk]) begin
          $fwrite(f, "Register (53,0) Value: %h\n", PRED53_0_buffer[clk]);
        end
        if (PRED53_1_buffer[clk] != PRED53_1_buffer[!clk]) begin
          $fwrite(f, "Register (53,1) Value: %h\n", PRED53_1_buffer[clk]);
        end
        if (PRED53_2_buffer[clk] != PRED53_2_buffer[!clk]) begin
          $fwrite(f, "Register (53,2) Value: %h\n", PRED53_2_buffer[clk]);
        end
        if (PRED53_3_buffer[clk] != PRED53_3_buffer[!clk]) begin
          $fwrite(f, "Register (53,3) Value: %h\n", PRED53_3_buffer[clk]);
        end
        if (PRED53_4_buffer[clk] != PRED53_4_buffer[!clk]) begin
          $fwrite(f, "Register (53,4) Value: %h\n", PRED53_4_buffer[clk]);
        end
        if (PRED53_5_buffer[clk] != PRED53_5_buffer[!clk]) begin
          $fwrite(f, "Register (53,5) Value: %h\n", PRED53_5_buffer[clk]);
        end
        if (PRED53_6_buffer[clk] != PRED53_6_buffer[!clk]) begin
          $fwrite(f, "Register (53,6) Value: %h\n", PRED53_6_buffer[clk]);
        end
        if (PRED53_7_buffer[clk] != PRED53_7_buffer[!clk]) begin
          $fwrite(f, "Register (53,7) Value: %h\n", PRED53_7_buffer[clk]);
        end
        if (PRED53_8_buffer[clk] != PRED53_8_buffer[!clk]) begin
          $fwrite(f, "Register (53,8) Value: %h\n", PRED53_8_buffer[clk]);
        end
        if (PRED53_9_buffer[clk] != PRED53_9_buffer[!clk]) begin
          $fwrite(f, "Register (53,9) Value: %h\n", PRED53_9_buffer[clk]);
        end
        if (PRED53_10_buffer[clk] != PRED53_10_buffer[!clk]) begin
          $fwrite(f, "Register (53,10) Value: %h\n", PRED53_10_buffer[clk]);
        end
        if (PRED53_11_buffer[clk] != PRED53_11_buffer[!clk]) begin
          $fwrite(f, "Register (53,11) Value: %h\n", PRED53_11_buffer[clk]);
        end
        if (PRED53_12_buffer[clk] != PRED53_12_buffer[!clk]) begin
          $fwrite(f, "Register (53,12) Value: %h\n", PRED53_12_buffer[clk]);
        end
        if (PRED53_13_buffer[clk] != PRED53_13_buffer[!clk]) begin
          $fwrite(f, "Register (53,13) Value: %h\n", PRED53_13_buffer[clk]);
        end
        if (PRED53_14_buffer[clk] != PRED53_14_buffer[!clk]) begin
          $fwrite(f, "Register (53,14) Value: %h\n", PRED53_14_buffer[clk]);
        end
        if (PRED53_15_buffer[clk] != PRED53_15_buffer[!clk]) begin
          $fwrite(f, "Register (53,15) Value: %h\n", PRED53_15_buffer[clk]);
        end
        if (PRED53_16_buffer[clk] != PRED53_16_buffer[!clk]) begin
          $fwrite(f, "Register (53,16) Value: %h\n", PRED53_16_buffer[clk]);
        end
        if (PRED53_17_buffer[clk] != PRED53_17_buffer[!clk]) begin
          $fwrite(f, "Register (53,17) Value: %h\n", PRED53_17_buffer[clk]);
        end
        if (PRED53_18_buffer[clk] != PRED53_18_buffer[!clk]) begin
          $fwrite(f, "Register (53,18) Value: %h\n", PRED53_18_buffer[clk]);
        end
        if (PRED53_19_buffer[clk] != PRED53_19_buffer[!clk]) begin
          $fwrite(f, "Register (53,19) Value: %h\n", PRED53_19_buffer[clk]);
        end
        if (PRED53_20_buffer[clk] != PRED53_20_buffer[!clk]) begin
          $fwrite(f, "Register (53,20) Value: %h\n", PRED53_20_buffer[clk]);
        end
        if (PRED53_21_buffer[clk] != PRED53_21_buffer[!clk]) begin
          $fwrite(f, "Register (53,21) Value: %h\n", PRED53_21_buffer[clk]);
        end
        if (PRED53_22_buffer[clk] != PRED53_22_buffer[!clk]) begin
          $fwrite(f, "Register (53,22) Value: %h\n", PRED53_22_buffer[clk]);
        end
        if (PRED53_23_buffer[clk] != PRED53_23_buffer[!clk]) begin
          $fwrite(f, "Register (53,23) Value: %h\n", PRED53_23_buffer[clk]);
        end
        if (PRED53_24_buffer[clk] != PRED53_24_buffer[!clk]) begin
          $fwrite(f, "Register (53,24) Value: %h\n", PRED53_24_buffer[clk]);
        end
        if (PRED53_25_buffer[clk] != PRED53_25_buffer[!clk]) begin
          $fwrite(f, "Register (53,25) Value: %h\n", PRED53_25_buffer[clk]);
        end
        if (PRED53_26_buffer[clk] != PRED53_26_buffer[!clk]) begin
          $fwrite(f, "Register (53,26) Value: %h\n", PRED53_26_buffer[clk]);
        end
        if (PRED53_27_buffer[clk] != PRED53_27_buffer[!clk]) begin
          $fwrite(f, "Register (53,27) Value: %h\n", PRED53_27_buffer[clk]);
        end
        if (PRED53_28_buffer[clk] != PRED53_28_buffer[!clk]) begin
          $fwrite(f, "Register (53,28) Value: %h\n", PRED53_28_buffer[clk]);
        end
        if (PRED53_29_buffer[clk] != PRED53_29_buffer[!clk]) begin
          $fwrite(f, "Register (53,29) Value: %h\n", PRED53_29_buffer[clk]);
        end
        if (PRED53_30_buffer[clk] != PRED53_30_buffer[!clk]) begin
          $fwrite(f, "Register (53,30) Value: %h\n", PRED53_30_buffer[clk]);
        end
        if (PRED53_31_buffer[clk] != PRED53_31_buffer[!clk]) begin
          $fwrite(f, "Register (53,31) Value: %h\n", PRED53_31_buffer[clk]);
        end
        if (PRED54_0_buffer[clk] != PRED54_0_buffer[!clk]) begin
          $fwrite(f, "Register (54,0) Value: %h\n", PRED54_0_buffer[clk]);
        end
        if (PRED54_1_buffer[clk] != PRED54_1_buffer[!clk]) begin
          $fwrite(f, "Register (54,1) Value: %h\n", PRED54_1_buffer[clk]);
        end
        if (PRED54_2_buffer[clk] != PRED54_2_buffer[!clk]) begin
          $fwrite(f, "Register (54,2) Value: %h\n", PRED54_2_buffer[clk]);
        end
        if (PRED54_3_buffer[clk] != PRED54_3_buffer[!clk]) begin
          $fwrite(f, "Register (54,3) Value: %h\n", PRED54_3_buffer[clk]);
        end
        if (PRED54_4_buffer[clk] != PRED54_4_buffer[!clk]) begin
          $fwrite(f, "Register (54,4) Value: %h\n", PRED54_4_buffer[clk]);
        end
        if (PRED54_5_buffer[clk] != PRED54_5_buffer[!clk]) begin
          $fwrite(f, "Register (54,5) Value: %h\n", PRED54_5_buffer[clk]);
        end
        if (PRED54_6_buffer[clk] != PRED54_6_buffer[!clk]) begin
          $fwrite(f, "Register (54,6) Value: %h\n", PRED54_6_buffer[clk]);
        end
        if (PRED54_7_buffer[clk] != PRED54_7_buffer[!clk]) begin
          $fwrite(f, "Register (54,7) Value: %h\n", PRED54_7_buffer[clk]);
        end
        if (PRED54_8_buffer[clk] != PRED54_8_buffer[!clk]) begin
          $fwrite(f, "Register (54,8) Value: %h\n", PRED54_8_buffer[clk]);
        end
        if (PRED54_9_buffer[clk] != PRED54_9_buffer[!clk]) begin
          $fwrite(f, "Register (54,9) Value: %h\n", PRED54_9_buffer[clk]);
        end
        if (PRED54_10_buffer[clk] != PRED54_10_buffer[!clk]) begin
          $fwrite(f, "Register (54,10) Value: %h\n", PRED54_10_buffer[clk]);
        end
        if (PRED54_11_buffer[clk] != PRED54_11_buffer[!clk]) begin
          $fwrite(f, "Register (54,11) Value: %h\n", PRED54_11_buffer[clk]);
        end
        if (PRED54_12_buffer[clk] != PRED54_12_buffer[!clk]) begin
          $fwrite(f, "Register (54,12) Value: %h\n", PRED54_12_buffer[clk]);
        end
        if (PRED54_13_buffer[clk] != PRED54_13_buffer[!clk]) begin
          $fwrite(f, "Register (54,13) Value: %h\n", PRED54_13_buffer[clk]);
        end
        if (PRED54_14_buffer[clk] != PRED54_14_buffer[!clk]) begin
          $fwrite(f, "Register (54,14) Value: %h\n", PRED54_14_buffer[clk]);
        end
        if (PRED54_15_buffer[clk] != PRED54_15_buffer[!clk]) begin
          $fwrite(f, "Register (54,15) Value: %h\n", PRED54_15_buffer[clk]);
        end
        if (PRED54_16_buffer[clk] != PRED54_16_buffer[!clk]) begin
          $fwrite(f, "Register (54,16) Value: %h\n", PRED54_16_buffer[clk]);
        end
        if (PRED54_17_buffer[clk] != PRED54_17_buffer[!clk]) begin
          $fwrite(f, "Register (54,17) Value: %h\n", PRED54_17_buffer[clk]);
        end
        if (PRED54_18_buffer[clk] != PRED54_18_buffer[!clk]) begin
          $fwrite(f, "Register (54,18) Value: %h\n", PRED54_18_buffer[clk]);
        end
        if (PRED54_19_buffer[clk] != PRED54_19_buffer[!clk]) begin
          $fwrite(f, "Register (54,19) Value: %h\n", PRED54_19_buffer[clk]);
        end
        if (PRED54_20_buffer[clk] != PRED54_20_buffer[!clk]) begin
          $fwrite(f, "Register (54,20) Value: %h\n", PRED54_20_buffer[clk]);
        end
        if (PRED54_21_buffer[clk] != PRED54_21_buffer[!clk]) begin
          $fwrite(f, "Register (54,21) Value: %h\n", PRED54_21_buffer[clk]);
        end
        if (PRED54_22_buffer[clk] != PRED54_22_buffer[!clk]) begin
          $fwrite(f, "Register (54,22) Value: %h\n", PRED54_22_buffer[clk]);
        end
        if (PRED54_23_buffer[clk] != PRED54_23_buffer[!clk]) begin
          $fwrite(f, "Register (54,23) Value: %h\n", PRED54_23_buffer[clk]);
        end
        if (PRED54_24_buffer[clk] != PRED54_24_buffer[!clk]) begin
          $fwrite(f, "Register (54,24) Value: %h\n", PRED54_24_buffer[clk]);
        end
        if (PRED54_25_buffer[clk] != PRED54_25_buffer[!clk]) begin
          $fwrite(f, "Register (54,25) Value: %h\n", PRED54_25_buffer[clk]);
        end
        if (PRED54_26_buffer[clk] != PRED54_26_buffer[!clk]) begin
          $fwrite(f, "Register (54,26) Value: %h\n", PRED54_26_buffer[clk]);
        end
        if (PRED54_27_buffer[clk] != PRED54_27_buffer[!clk]) begin
          $fwrite(f, "Register (54,27) Value: %h\n", PRED54_27_buffer[clk]);
        end
        if (PRED54_28_buffer[clk] != PRED54_28_buffer[!clk]) begin
          $fwrite(f, "Register (54,28) Value: %h\n", PRED54_28_buffer[clk]);
        end
        if (PRED54_29_buffer[clk] != PRED54_29_buffer[!clk]) begin
          $fwrite(f, "Register (54,29) Value: %h\n", PRED54_29_buffer[clk]);
        end
        if (PRED54_30_buffer[clk] != PRED54_30_buffer[!clk]) begin
          $fwrite(f, "Register (54,30) Value: %h\n", PRED54_30_buffer[clk]);
        end
        if (PRED54_31_buffer[clk] != PRED54_31_buffer[!clk]) begin
          $fwrite(f, "Register (54,31) Value: %h\n", PRED54_31_buffer[clk]);
        end
        if (PRED55_0_buffer[clk] != PRED55_0_buffer[!clk]) begin
          $fwrite(f, "Register (55,0) Value: %h\n", PRED55_0_buffer[clk]);
        end
        if (PRED55_1_buffer[clk] != PRED55_1_buffer[!clk]) begin
          $fwrite(f, "Register (55,1) Value: %h\n", PRED55_1_buffer[clk]);
        end
        if (PRED55_2_buffer[clk] != PRED55_2_buffer[!clk]) begin
          $fwrite(f, "Register (55,2) Value: %h\n", PRED55_2_buffer[clk]);
        end
        if (PRED55_3_buffer[clk] != PRED55_3_buffer[!clk]) begin
          $fwrite(f, "Register (55,3) Value: %h\n", PRED55_3_buffer[clk]);
        end
        if (PRED55_4_buffer[clk] != PRED55_4_buffer[!clk]) begin
          $fwrite(f, "Register (55,4) Value: %h\n", PRED55_4_buffer[clk]);
        end
        if (PRED55_5_buffer[clk] != PRED55_5_buffer[!clk]) begin
          $fwrite(f, "Register (55,5) Value: %h\n", PRED55_5_buffer[clk]);
        end
        if (PRED55_6_buffer[clk] != PRED55_6_buffer[!clk]) begin
          $fwrite(f, "Register (55,6) Value: %h\n", PRED55_6_buffer[clk]);
        end
        if (PRED55_7_buffer[clk] != PRED55_7_buffer[!clk]) begin
          $fwrite(f, "Register (55,7) Value: %h\n", PRED55_7_buffer[clk]);
        end
        if (PRED55_8_buffer[clk] != PRED55_8_buffer[!clk]) begin
          $fwrite(f, "Register (55,8) Value: %h\n", PRED55_8_buffer[clk]);
        end
        if (PRED55_9_buffer[clk] != PRED55_9_buffer[!clk]) begin
          $fwrite(f, "Register (55,9) Value: %h\n", PRED55_9_buffer[clk]);
        end
        if (PRED55_10_buffer[clk] != PRED55_10_buffer[!clk]) begin
          $fwrite(f, "Register (55,10) Value: %h\n", PRED55_10_buffer[clk]);
        end
        if (PRED55_11_buffer[clk] != PRED55_11_buffer[!clk]) begin
          $fwrite(f, "Register (55,11) Value: %h\n", PRED55_11_buffer[clk]);
        end
        if (PRED55_12_buffer[clk] != PRED55_12_buffer[!clk]) begin
          $fwrite(f, "Register (55,12) Value: %h\n", PRED55_12_buffer[clk]);
        end
        if (PRED55_13_buffer[clk] != PRED55_13_buffer[!clk]) begin
          $fwrite(f, "Register (55,13) Value: %h\n", PRED55_13_buffer[clk]);
        end
        if (PRED55_14_buffer[clk] != PRED55_14_buffer[!clk]) begin
          $fwrite(f, "Register (55,14) Value: %h\n", PRED55_14_buffer[clk]);
        end
        if (PRED55_15_buffer[clk] != PRED55_15_buffer[!clk]) begin
          $fwrite(f, "Register (55,15) Value: %h\n", PRED55_15_buffer[clk]);
        end
        if (PRED55_16_buffer[clk] != PRED55_16_buffer[!clk]) begin
          $fwrite(f, "Register (55,16) Value: %h\n", PRED55_16_buffer[clk]);
        end
        if (PRED55_17_buffer[clk] != PRED55_17_buffer[!clk]) begin
          $fwrite(f, "Register (55,17) Value: %h\n", PRED55_17_buffer[clk]);
        end
        if (PRED55_18_buffer[clk] != PRED55_18_buffer[!clk]) begin
          $fwrite(f, "Register (55,18) Value: %h\n", PRED55_18_buffer[clk]);
        end
        if (PRED55_19_buffer[clk] != PRED55_19_buffer[!clk]) begin
          $fwrite(f, "Register (55,19) Value: %h\n", PRED55_19_buffer[clk]);
        end
        if (PRED55_20_buffer[clk] != PRED55_20_buffer[!clk]) begin
          $fwrite(f, "Register (55,20) Value: %h\n", PRED55_20_buffer[clk]);
        end
        if (PRED55_21_buffer[clk] != PRED55_21_buffer[!clk]) begin
          $fwrite(f, "Register (55,21) Value: %h\n", PRED55_21_buffer[clk]);
        end
        if (PRED55_22_buffer[clk] != PRED55_22_buffer[!clk]) begin
          $fwrite(f, "Register (55,22) Value: %h\n", PRED55_22_buffer[clk]);
        end
        if (PRED55_23_buffer[clk] != PRED55_23_buffer[!clk]) begin
          $fwrite(f, "Register (55,23) Value: %h\n", PRED55_23_buffer[clk]);
        end
        if (PRED55_24_buffer[clk] != PRED55_24_buffer[!clk]) begin
          $fwrite(f, "Register (55,24) Value: %h\n", PRED55_24_buffer[clk]);
        end
        if (PRED55_25_buffer[clk] != PRED55_25_buffer[!clk]) begin
          $fwrite(f, "Register (55,25) Value: %h\n", PRED55_25_buffer[clk]);
        end
        if (PRED55_26_buffer[clk] != PRED55_26_buffer[!clk]) begin
          $fwrite(f, "Register (55,26) Value: %h\n", PRED55_26_buffer[clk]);
        end
        if (PRED55_27_buffer[clk] != PRED55_27_buffer[!clk]) begin
          $fwrite(f, "Register (55,27) Value: %h\n", PRED55_27_buffer[clk]);
        end
        if (PRED55_28_buffer[clk] != PRED55_28_buffer[!clk]) begin
          $fwrite(f, "Register (55,28) Value: %h\n", PRED55_28_buffer[clk]);
        end
        if (PRED55_29_buffer[clk] != PRED55_29_buffer[!clk]) begin
          $fwrite(f, "Register (55,29) Value: %h\n", PRED55_29_buffer[clk]);
        end
        if (PRED55_30_buffer[clk] != PRED55_30_buffer[!clk]) begin
          $fwrite(f, "Register (55,30) Value: %h\n", PRED55_30_buffer[clk]);
        end
        if (PRED55_31_buffer[clk] != PRED55_31_buffer[!clk]) begin
          $fwrite(f, "Register (55,31) Value: %h\n", PRED55_31_buffer[clk]);
        end
        if (PRED56_0_buffer[clk] != PRED56_0_buffer[!clk]) begin
          $fwrite(f, "Register (56,0) Value: %h\n", PRED56_0_buffer[clk]);
        end
        if (PRED56_1_buffer[clk] != PRED56_1_buffer[!clk]) begin
          $fwrite(f, "Register (56,1) Value: %h\n", PRED56_1_buffer[clk]);
        end
        if (PRED56_2_buffer[clk] != PRED56_2_buffer[!clk]) begin
          $fwrite(f, "Register (56,2) Value: %h\n", PRED56_2_buffer[clk]);
        end
        if (PRED56_3_buffer[clk] != PRED56_3_buffer[!clk]) begin
          $fwrite(f, "Register (56,3) Value: %h\n", PRED56_3_buffer[clk]);
        end
        if (PRED56_4_buffer[clk] != PRED56_4_buffer[!clk]) begin
          $fwrite(f, "Register (56,4) Value: %h\n", PRED56_4_buffer[clk]);
        end
        if (PRED56_5_buffer[clk] != PRED56_5_buffer[!clk]) begin
          $fwrite(f, "Register (56,5) Value: %h\n", PRED56_5_buffer[clk]);
        end
        if (PRED56_6_buffer[clk] != PRED56_6_buffer[!clk]) begin
          $fwrite(f, "Register (56,6) Value: %h\n", PRED56_6_buffer[clk]);
        end
        if (PRED56_7_buffer[clk] != PRED56_7_buffer[!clk]) begin
          $fwrite(f, "Register (56,7) Value: %h\n", PRED56_7_buffer[clk]);
        end
        if (PRED56_8_buffer[clk] != PRED56_8_buffer[!clk]) begin
          $fwrite(f, "Register (56,8) Value: %h\n", PRED56_8_buffer[clk]);
        end
        if (PRED56_9_buffer[clk] != PRED56_9_buffer[!clk]) begin
          $fwrite(f, "Register (56,9) Value: %h\n", PRED56_9_buffer[clk]);
        end
        if (PRED56_10_buffer[clk] != PRED56_10_buffer[!clk]) begin
          $fwrite(f, "Register (56,10) Value: %h\n", PRED56_10_buffer[clk]);
        end
        if (PRED56_11_buffer[clk] != PRED56_11_buffer[!clk]) begin
          $fwrite(f, "Register (56,11) Value: %h\n", PRED56_11_buffer[clk]);
        end
        if (PRED56_12_buffer[clk] != PRED56_12_buffer[!clk]) begin
          $fwrite(f, "Register (56,12) Value: %h\n", PRED56_12_buffer[clk]);
        end
        if (PRED56_13_buffer[clk] != PRED56_13_buffer[!clk]) begin
          $fwrite(f, "Register (56,13) Value: %h\n", PRED56_13_buffer[clk]);
        end
        if (PRED56_14_buffer[clk] != PRED56_14_buffer[!clk]) begin
          $fwrite(f, "Register (56,14) Value: %h\n", PRED56_14_buffer[clk]);
        end
        if (PRED56_15_buffer[clk] != PRED56_15_buffer[!clk]) begin
          $fwrite(f, "Register (56,15) Value: %h\n", PRED56_15_buffer[clk]);
        end
        if (PRED56_16_buffer[clk] != PRED56_16_buffer[!clk]) begin
          $fwrite(f, "Register (56,16) Value: %h\n", PRED56_16_buffer[clk]);
        end
        if (PRED56_17_buffer[clk] != PRED56_17_buffer[!clk]) begin
          $fwrite(f, "Register (56,17) Value: %h\n", PRED56_17_buffer[clk]);
        end
        if (PRED56_18_buffer[clk] != PRED56_18_buffer[!clk]) begin
          $fwrite(f, "Register (56,18) Value: %h\n", PRED56_18_buffer[clk]);
        end
        if (PRED56_19_buffer[clk] != PRED56_19_buffer[!clk]) begin
          $fwrite(f, "Register (56,19) Value: %h\n", PRED56_19_buffer[clk]);
        end
        if (PRED56_20_buffer[clk] != PRED56_20_buffer[!clk]) begin
          $fwrite(f, "Register (56,20) Value: %h\n", PRED56_20_buffer[clk]);
        end
        if (PRED56_21_buffer[clk] != PRED56_21_buffer[!clk]) begin
          $fwrite(f, "Register (56,21) Value: %h\n", PRED56_21_buffer[clk]);
        end
        if (PRED56_22_buffer[clk] != PRED56_22_buffer[!clk]) begin
          $fwrite(f, "Register (56,22) Value: %h\n", PRED56_22_buffer[clk]);
        end
        if (PRED56_23_buffer[clk] != PRED56_23_buffer[!clk]) begin
          $fwrite(f, "Register (56,23) Value: %h\n", PRED56_23_buffer[clk]);
        end
        if (PRED56_24_buffer[clk] != PRED56_24_buffer[!clk]) begin
          $fwrite(f, "Register (56,24) Value: %h\n", PRED56_24_buffer[clk]);
        end
        if (PRED56_25_buffer[clk] != PRED56_25_buffer[!clk]) begin
          $fwrite(f, "Register (56,25) Value: %h\n", PRED56_25_buffer[clk]);
        end
        if (PRED56_26_buffer[clk] != PRED56_26_buffer[!clk]) begin
          $fwrite(f, "Register (56,26) Value: %h\n", PRED56_26_buffer[clk]);
        end
        if (PRED56_27_buffer[clk] != PRED56_27_buffer[!clk]) begin
          $fwrite(f, "Register (56,27) Value: %h\n", PRED56_27_buffer[clk]);
        end
        if (PRED56_28_buffer[clk] != PRED56_28_buffer[!clk]) begin
          $fwrite(f, "Register (56,28) Value: %h\n", PRED56_28_buffer[clk]);
        end
        if (PRED56_29_buffer[clk] != PRED56_29_buffer[!clk]) begin
          $fwrite(f, "Register (56,29) Value: %h\n", PRED56_29_buffer[clk]);
        end
        if (PRED56_30_buffer[clk] != PRED56_30_buffer[!clk]) begin
          $fwrite(f, "Register (56,30) Value: %h\n", PRED56_30_buffer[clk]);
        end
        if (PRED56_31_buffer[clk] != PRED56_31_buffer[!clk]) begin
          $fwrite(f, "Register (56,31) Value: %h\n", PRED56_31_buffer[clk]);
        end
        if (PRED57_0_buffer[clk] != PRED57_0_buffer[!clk]) begin
          $fwrite(f, "Register (57,0) Value: %h\n", PRED57_0_buffer[clk]);
        end
        if (PRED57_1_buffer[clk] != PRED57_1_buffer[!clk]) begin
          $fwrite(f, "Register (57,1) Value: %h\n", PRED57_1_buffer[clk]);
        end
        if (PRED57_2_buffer[clk] != PRED57_2_buffer[!clk]) begin
          $fwrite(f, "Register (57,2) Value: %h\n", PRED57_2_buffer[clk]);
        end
        if (PRED57_3_buffer[clk] != PRED57_3_buffer[!clk]) begin
          $fwrite(f, "Register (57,3) Value: %h\n", PRED57_3_buffer[clk]);
        end
        if (PRED57_4_buffer[clk] != PRED57_4_buffer[!clk]) begin
          $fwrite(f, "Register (57,4) Value: %h\n", PRED57_4_buffer[clk]);
        end
        if (PRED57_5_buffer[clk] != PRED57_5_buffer[!clk]) begin
          $fwrite(f, "Register (57,5) Value: %h\n", PRED57_5_buffer[clk]);
        end
        if (PRED57_6_buffer[clk] != PRED57_6_buffer[!clk]) begin
          $fwrite(f, "Register (57,6) Value: %h\n", PRED57_6_buffer[clk]);
        end
        if (PRED57_7_buffer[clk] != PRED57_7_buffer[!clk]) begin
          $fwrite(f, "Register (57,7) Value: %h\n", PRED57_7_buffer[clk]);
        end
        if (PRED57_8_buffer[clk] != PRED57_8_buffer[!clk]) begin
          $fwrite(f, "Register (57,8) Value: %h\n", PRED57_8_buffer[clk]);
        end
        if (PRED57_9_buffer[clk] != PRED57_9_buffer[!clk]) begin
          $fwrite(f, "Register (57,9) Value: %h\n", PRED57_9_buffer[clk]);
        end
        if (PRED57_10_buffer[clk] != PRED57_10_buffer[!clk]) begin
          $fwrite(f, "Register (57,10) Value: %h\n", PRED57_10_buffer[clk]);
        end
        if (PRED57_11_buffer[clk] != PRED57_11_buffer[!clk]) begin
          $fwrite(f, "Register (57,11) Value: %h\n", PRED57_11_buffer[clk]);
        end
        if (PRED57_12_buffer[clk] != PRED57_12_buffer[!clk]) begin
          $fwrite(f, "Register (57,12) Value: %h\n", PRED57_12_buffer[clk]);
        end
        if (PRED57_13_buffer[clk] != PRED57_13_buffer[!clk]) begin
          $fwrite(f, "Register (57,13) Value: %h\n", PRED57_13_buffer[clk]);
        end
        if (PRED57_14_buffer[clk] != PRED57_14_buffer[!clk]) begin
          $fwrite(f, "Register (57,14) Value: %h\n", PRED57_14_buffer[clk]);
        end
        if (PRED57_15_buffer[clk] != PRED57_15_buffer[!clk]) begin
          $fwrite(f, "Register (57,15) Value: %h\n", PRED57_15_buffer[clk]);
        end
        if (PRED57_16_buffer[clk] != PRED57_16_buffer[!clk]) begin
          $fwrite(f, "Register (57,16) Value: %h\n", PRED57_16_buffer[clk]);
        end
        if (PRED57_17_buffer[clk] != PRED57_17_buffer[!clk]) begin
          $fwrite(f, "Register (57,17) Value: %h\n", PRED57_17_buffer[clk]);
        end
        if (PRED57_18_buffer[clk] != PRED57_18_buffer[!clk]) begin
          $fwrite(f, "Register (57,18) Value: %h\n", PRED57_18_buffer[clk]);
        end
        if (PRED57_19_buffer[clk] != PRED57_19_buffer[!clk]) begin
          $fwrite(f, "Register (57,19) Value: %h\n", PRED57_19_buffer[clk]);
        end
        if (PRED57_20_buffer[clk] != PRED57_20_buffer[!clk]) begin
          $fwrite(f, "Register (57,20) Value: %h\n", PRED57_20_buffer[clk]);
        end
        if (PRED57_21_buffer[clk] != PRED57_21_buffer[!clk]) begin
          $fwrite(f, "Register (57,21) Value: %h\n", PRED57_21_buffer[clk]);
        end
        if (PRED57_22_buffer[clk] != PRED57_22_buffer[!clk]) begin
          $fwrite(f, "Register (57,22) Value: %h\n", PRED57_22_buffer[clk]);
        end
        if (PRED57_23_buffer[clk] != PRED57_23_buffer[!clk]) begin
          $fwrite(f, "Register (57,23) Value: %h\n", PRED57_23_buffer[clk]);
        end
        if (PRED57_24_buffer[clk] != PRED57_24_buffer[!clk]) begin
          $fwrite(f, "Register (57,24) Value: %h\n", PRED57_24_buffer[clk]);
        end
        if (PRED57_25_buffer[clk] != PRED57_25_buffer[!clk]) begin
          $fwrite(f, "Register (57,25) Value: %h\n", PRED57_25_buffer[clk]);
        end
        if (PRED57_26_buffer[clk] != PRED57_26_buffer[!clk]) begin
          $fwrite(f, "Register (57,26) Value: %h\n", PRED57_26_buffer[clk]);
        end
        if (PRED57_27_buffer[clk] != PRED57_27_buffer[!clk]) begin
          $fwrite(f, "Register (57,27) Value: %h\n", PRED57_27_buffer[clk]);
        end
        if (PRED57_28_buffer[clk] != PRED57_28_buffer[!clk]) begin
          $fwrite(f, "Register (57,28) Value: %h\n", PRED57_28_buffer[clk]);
        end
        if (PRED57_29_buffer[clk] != PRED57_29_buffer[!clk]) begin
          $fwrite(f, "Register (57,29) Value: %h\n", PRED57_29_buffer[clk]);
        end
        if (PRED57_30_buffer[clk] != PRED57_30_buffer[!clk]) begin
          $fwrite(f, "Register (57,30) Value: %h\n", PRED57_30_buffer[clk]);
        end
        if (PRED57_31_buffer[clk] != PRED57_31_buffer[!clk]) begin
          $fwrite(f, "Register (57,31) Value: %h\n", PRED57_31_buffer[clk]);
        end
        if (PRED58_0_buffer[clk] != PRED58_0_buffer[!clk]) begin
          $fwrite(f, "Register (58,0) Value: %h\n", PRED58_0_buffer[clk]);
        end
        if (PRED58_1_buffer[clk] != PRED58_1_buffer[!clk]) begin
          $fwrite(f, "Register (58,1) Value: %h\n", PRED58_1_buffer[clk]);
        end
        if (PRED58_2_buffer[clk] != PRED58_2_buffer[!clk]) begin
          $fwrite(f, "Register (58,2) Value: %h\n", PRED58_2_buffer[clk]);
        end
        if (PRED58_3_buffer[clk] != PRED58_3_buffer[!clk]) begin
          $fwrite(f, "Register (58,3) Value: %h\n", PRED58_3_buffer[clk]);
        end
        if (PRED58_4_buffer[clk] != PRED58_4_buffer[!clk]) begin
          $fwrite(f, "Register (58,4) Value: %h\n", PRED58_4_buffer[clk]);
        end
        if (PRED58_5_buffer[clk] != PRED58_5_buffer[!clk]) begin
          $fwrite(f, "Register (58,5) Value: %h\n", PRED58_5_buffer[clk]);
        end
        if (PRED58_6_buffer[clk] != PRED58_6_buffer[!clk]) begin
          $fwrite(f, "Register (58,6) Value: %h\n", PRED58_6_buffer[clk]);
        end
        if (PRED58_7_buffer[clk] != PRED58_7_buffer[!clk]) begin
          $fwrite(f, "Register (58,7) Value: %h\n", PRED58_7_buffer[clk]);
        end
        if (PRED58_8_buffer[clk] != PRED58_8_buffer[!clk]) begin
          $fwrite(f, "Register (58,8) Value: %h\n", PRED58_8_buffer[clk]);
        end
        if (PRED58_9_buffer[clk] != PRED58_9_buffer[!clk]) begin
          $fwrite(f, "Register (58,9) Value: %h\n", PRED58_9_buffer[clk]);
        end
        if (PRED58_10_buffer[clk] != PRED58_10_buffer[!clk]) begin
          $fwrite(f, "Register (58,10) Value: %h\n", PRED58_10_buffer[clk]);
        end
        if (PRED58_11_buffer[clk] != PRED58_11_buffer[!clk]) begin
          $fwrite(f, "Register (58,11) Value: %h\n", PRED58_11_buffer[clk]);
        end
        if (PRED58_12_buffer[clk] != PRED58_12_buffer[!clk]) begin
          $fwrite(f, "Register (58,12) Value: %h\n", PRED58_12_buffer[clk]);
        end
        if (PRED58_13_buffer[clk] != PRED58_13_buffer[!clk]) begin
          $fwrite(f, "Register (58,13) Value: %h\n", PRED58_13_buffer[clk]);
        end
        if (PRED58_14_buffer[clk] != PRED58_14_buffer[!clk]) begin
          $fwrite(f, "Register (58,14) Value: %h\n", PRED58_14_buffer[clk]);
        end
        if (PRED58_15_buffer[clk] != PRED58_15_buffer[!clk]) begin
          $fwrite(f, "Register (58,15) Value: %h\n", PRED58_15_buffer[clk]);
        end
        if (PRED58_16_buffer[clk] != PRED58_16_buffer[!clk]) begin
          $fwrite(f, "Register (58,16) Value: %h\n", PRED58_16_buffer[clk]);
        end
        if (PRED58_17_buffer[clk] != PRED58_17_buffer[!clk]) begin
          $fwrite(f, "Register (58,17) Value: %h\n", PRED58_17_buffer[clk]);
        end
        if (PRED58_18_buffer[clk] != PRED58_18_buffer[!clk]) begin
          $fwrite(f, "Register (58,18) Value: %h\n", PRED58_18_buffer[clk]);
        end
        if (PRED58_19_buffer[clk] != PRED58_19_buffer[!clk]) begin
          $fwrite(f, "Register (58,19) Value: %h\n", PRED58_19_buffer[clk]);
        end
        if (PRED58_20_buffer[clk] != PRED58_20_buffer[!clk]) begin
          $fwrite(f, "Register (58,20) Value: %h\n", PRED58_20_buffer[clk]);
        end
        if (PRED58_21_buffer[clk] != PRED58_21_buffer[!clk]) begin
          $fwrite(f, "Register (58,21) Value: %h\n", PRED58_21_buffer[clk]);
        end
        if (PRED58_22_buffer[clk] != PRED58_22_buffer[!clk]) begin
          $fwrite(f, "Register (58,22) Value: %h\n", PRED58_22_buffer[clk]);
        end
        if (PRED58_23_buffer[clk] != PRED58_23_buffer[!clk]) begin
          $fwrite(f, "Register (58,23) Value: %h\n", PRED58_23_buffer[clk]);
        end
        if (PRED58_24_buffer[clk] != PRED58_24_buffer[!clk]) begin
          $fwrite(f, "Register (58,24) Value: %h\n", PRED58_24_buffer[clk]);
        end
        if (PRED58_25_buffer[clk] != PRED58_25_buffer[!clk]) begin
          $fwrite(f, "Register (58,25) Value: %h\n", PRED58_25_buffer[clk]);
        end
        if (PRED58_26_buffer[clk] != PRED58_26_buffer[!clk]) begin
          $fwrite(f, "Register (58,26) Value: %h\n", PRED58_26_buffer[clk]);
        end
        if (PRED58_27_buffer[clk] != PRED58_27_buffer[!clk]) begin
          $fwrite(f, "Register (58,27) Value: %h\n", PRED58_27_buffer[clk]);
        end
        if (PRED58_28_buffer[clk] != PRED58_28_buffer[!clk]) begin
          $fwrite(f, "Register (58,28) Value: %h\n", PRED58_28_buffer[clk]);
        end
        if (PRED58_29_buffer[clk] != PRED58_29_buffer[!clk]) begin
          $fwrite(f, "Register (58,29) Value: %h\n", PRED58_29_buffer[clk]);
        end
        if (PRED58_30_buffer[clk] != PRED58_30_buffer[!clk]) begin
          $fwrite(f, "Register (58,30) Value: %h\n", PRED58_30_buffer[clk]);
        end
        if (PRED58_31_buffer[clk] != PRED58_31_buffer[!clk]) begin
          $fwrite(f, "Register (58,31) Value: %h\n", PRED58_31_buffer[clk]);
        end
        if (PRED59_0_buffer[clk] != PRED59_0_buffer[!clk]) begin
          $fwrite(f, "Register (59,0) Value: %h\n", PRED59_0_buffer[clk]);
        end
        if (PRED59_1_buffer[clk] != PRED59_1_buffer[!clk]) begin
          $fwrite(f, "Register (59,1) Value: %h\n", PRED59_1_buffer[clk]);
        end
        if (PRED59_2_buffer[clk] != PRED59_2_buffer[!clk]) begin
          $fwrite(f, "Register (59,2) Value: %h\n", PRED59_2_buffer[clk]);
        end
        if (PRED59_3_buffer[clk] != PRED59_3_buffer[!clk]) begin
          $fwrite(f, "Register (59,3) Value: %h\n", PRED59_3_buffer[clk]);
        end
        if (PRED59_4_buffer[clk] != PRED59_4_buffer[!clk]) begin
          $fwrite(f, "Register (59,4) Value: %h\n", PRED59_4_buffer[clk]);
        end
        if (PRED59_5_buffer[clk] != PRED59_5_buffer[!clk]) begin
          $fwrite(f, "Register (59,5) Value: %h\n", PRED59_5_buffer[clk]);
        end
        if (PRED59_6_buffer[clk] != PRED59_6_buffer[!clk]) begin
          $fwrite(f, "Register (59,6) Value: %h\n", PRED59_6_buffer[clk]);
        end
        if (PRED59_7_buffer[clk] != PRED59_7_buffer[!clk]) begin
          $fwrite(f, "Register (59,7) Value: %h\n", PRED59_7_buffer[clk]);
        end
        if (PRED59_8_buffer[clk] != PRED59_8_buffer[!clk]) begin
          $fwrite(f, "Register (59,8) Value: %h\n", PRED59_8_buffer[clk]);
        end
        if (PRED59_9_buffer[clk] != PRED59_9_buffer[!clk]) begin
          $fwrite(f, "Register (59,9) Value: %h\n", PRED59_9_buffer[clk]);
        end
        if (PRED59_10_buffer[clk] != PRED59_10_buffer[!clk]) begin
          $fwrite(f, "Register (59,10) Value: %h\n", PRED59_10_buffer[clk]);
        end
        if (PRED59_11_buffer[clk] != PRED59_11_buffer[!clk]) begin
          $fwrite(f, "Register (59,11) Value: %h\n", PRED59_11_buffer[clk]);
        end
        if (PRED59_12_buffer[clk] != PRED59_12_buffer[!clk]) begin
          $fwrite(f, "Register (59,12) Value: %h\n", PRED59_12_buffer[clk]);
        end
        if (PRED59_13_buffer[clk] != PRED59_13_buffer[!clk]) begin
          $fwrite(f, "Register (59,13) Value: %h\n", PRED59_13_buffer[clk]);
        end
        if (PRED59_14_buffer[clk] != PRED59_14_buffer[!clk]) begin
          $fwrite(f, "Register (59,14) Value: %h\n", PRED59_14_buffer[clk]);
        end
        if (PRED59_15_buffer[clk] != PRED59_15_buffer[!clk]) begin
          $fwrite(f, "Register (59,15) Value: %h\n", PRED59_15_buffer[clk]);
        end
        if (PRED59_16_buffer[clk] != PRED59_16_buffer[!clk]) begin
          $fwrite(f, "Register (59,16) Value: %h\n", PRED59_16_buffer[clk]);
        end
        if (PRED59_17_buffer[clk] != PRED59_17_buffer[!clk]) begin
          $fwrite(f, "Register (59,17) Value: %h\n", PRED59_17_buffer[clk]);
        end
        if (PRED59_18_buffer[clk] != PRED59_18_buffer[!clk]) begin
          $fwrite(f, "Register (59,18) Value: %h\n", PRED59_18_buffer[clk]);
        end
        if (PRED59_19_buffer[clk] != PRED59_19_buffer[!clk]) begin
          $fwrite(f, "Register (59,19) Value: %h\n", PRED59_19_buffer[clk]);
        end
        if (PRED59_20_buffer[clk] != PRED59_20_buffer[!clk]) begin
          $fwrite(f, "Register (59,20) Value: %h\n", PRED59_20_buffer[clk]);
        end
        if (PRED59_21_buffer[clk] != PRED59_21_buffer[!clk]) begin
          $fwrite(f, "Register (59,21) Value: %h\n", PRED59_21_buffer[clk]);
        end
        if (PRED59_22_buffer[clk] != PRED59_22_buffer[!clk]) begin
          $fwrite(f, "Register (59,22) Value: %h\n", PRED59_22_buffer[clk]);
        end
        if (PRED59_23_buffer[clk] != PRED59_23_buffer[!clk]) begin
          $fwrite(f, "Register (59,23) Value: %h\n", PRED59_23_buffer[clk]);
        end
        if (PRED59_24_buffer[clk] != PRED59_24_buffer[!clk]) begin
          $fwrite(f, "Register (59,24) Value: %h\n", PRED59_24_buffer[clk]);
        end
        if (PRED59_25_buffer[clk] != PRED59_25_buffer[!clk]) begin
          $fwrite(f, "Register (59,25) Value: %h\n", PRED59_25_buffer[clk]);
        end
        if (PRED59_26_buffer[clk] != PRED59_26_buffer[!clk]) begin
          $fwrite(f, "Register (59,26) Value: %h\n", PRED59_26_buffer[clk]);
        end
        if (PRED59_27_buffer[clk] != PRED59_27_buffer[!clk]) begin
          $fwrite(f, "Register (59,27) Value: %h\n", PRED59_27_buffer[clk]);
        end
        if (PRED59_28_buffer[clk] != PRED59_28_buffer[!clk]) begin
          $fwrite(f, "Register (59,28) Value: %h\n", PRED59_28_buffer[clk]);
        end
        if (PRED59_29_buffer[clk] != PRED59_29_buffer[!clk]) begin
          $fwrite(f, "Register (59,29) Value: %h\n", PRED59_29_buffer[clk]);
        end
        if (PRED59_30_buffer[clk] != PRED59_30_buffer[!clk]) begin
          $fwrite(f, "Register (59,30) Value: %h\n", PRED59_30_buffer[clk]);
        end
        if (PRED59_31_buffer[clk] != PRED59_31_buffer[!clk]) begin
          $fwrite(f, "Register (59,31) Value: %h\n", PRED59_31_buffer[clk]);
        end
        if (PRED60_0_buffer[clk] != PRED60_0_buffer[!clk]) begin
          $fwrite(f, "Register (60,0) Value: %h\n", PRED60_0_buffer[clk]);
        end
        if (PRED60_1_buffer[clk] != PRED60_1_buffer[!clk]) begin
          $fwrite(f, "Register (60,1) Value: %h\n", PRED60_1_buffer[clk]);
        end
        if (PRED60_2_buffer[clk] != PRED60_2_buffer[!clk]) begin
          $fwrite(f, "Register (60,2) Value: %h\n", PRED60_2_buffer[clk]);
        end
        if (PRED60_3_buffer[clk] != PRED60_3_buffer[!clk]) begin
          $fwrite(f, "Register (60,3) Value: %h\n", PRED60_3_buffer[clk]);
        end
        if (PRED60_4_buffer[clk] != PRED60_4_buffer[!clk]) begin
          $fwrite(f, "Register (60,4) Value: %h\n", PRED60_4_buffer[clk]);
        end
        if (PRED60_5_buffer[clk] != PRED60_5_buffer[!clk]) begin
          $fwrite(f, "Register (60,5) Value: %h\n", PRED60_5_buffer[clk]);
        end
        if (PRED60_6_buffer[clk] != PRED60_6_buffer[!clk]) begin
          $fwrite(f, "Register (60,6) Value: %h\n", PRED60_6_buffer[clk]);
        end
        if (PRED60_7_buffer[clk] != PRED60_7_buffer[!clk]) begin
          $fwrite(f, "Register (60,7) Value: %h\n", PRED60_7_buffer[clk]);
        end
        if (PRED60_8_buffer[clk] != PRED60_8_buffer[!clk]) begin
          $fwrite(f, "Register (60,8) Value: %h\n", PRED60_8_buffer[clk]);
        end
        if (PRED60_9_buffer[clk] != PRED60_9_buffer[!clk]) begin
          $fwrite(f, "Register (60,9) Value: %h\n", PRED60_9_buffer[clk]);
        end
        if (PRED60_10_buffer[clk] != PRED60_10_buffer[!clk]) begin
          $fwrite(f, "Register (60,10) Value: %h\n", PRED60_10_buffer[clk]);
        end
        if (PRED60_11_buffer[clk] != PRED60_11_buffer[!clk]) begin
          $fwrite(f, "Register (60,11) Value: %h\n", PRED60_11_buffer[clk]);
        end
        if (PRED60_12_buffer[clk] != PRED60_12_buffer[!clk]) begin
          $fwrite(f, "Register (60,12) Value: %h\n", PRED60_12_buffer[clk]);
        end
        if (PRED60_13_buffer[clk] != PRED60_13_buffer[!clk]) begin
          $fwrite(f, "Register (60,13) Value: %h\n", PRED60_13_buffer[clk]);
        end
        if (PRED60_14_buffer[clk] != PRED60_14_buffer[!clk]) begin
          $fwrite(f, "Register (60,14) Value: %h\n", PRED60_14_buffer[clk]);
        end
        if (PRED60_15_buffer[clk] != PRED60_15_buffer[!clk]) begin
          $fwrite(f, "Register (60,15) Value: %h\n", PRED60_15_buffer[clk]);
        end
        if (PRED60_16_buffer[clk] != PRED60_16_buffer[!clk]) begin
          $fwrite(f, "Register (60,16) Value: %h\n", PRED60_16_buffer[clk]);
        end
        if (PRED60_17_buffer[clk] != PRED60_17_buffer[!clk]) begin
          $fwrite(f, "Register (60,17) Value: %h\n", PRED60_17_buffer[clk]);
        end
        if (PRED60_18_buffer[clk] != PRED60_18_buffer[!clk]) begin
          $fwrite(f, "Register (60,18) Value: %h\n", PRED60_18_buffer[clk]);
        end
        if (PRED60_19_buffer[clk] != PRED60_19_buffer[!clk]) begin
          $fwrite(f, "Register (60,19) Value: %h\n", PRED60_19_buffer[clk]);
        end
        if (PRED60_20_buffer[clk] != PRED60_20_buffer[!clk]) begin
          $fwrite(f, "Register (60,20) Value: %h\n", PRED60_20_buffer[clk]);
        end
        if (PRED60_21_buffer[clk] != PRED60_21_buffer[!clk]) begin
          $fwrite(f, "Register (60,21) Value: %h\n", PRED60_21_buffer[clk]);
        end
        if (PRED60_22_buffer[clk] != PRED60_22_buffer[!clk]) begin
          $fwrite(f, "Register (60,22) Value: %h\n", PRED60_22_buffer[clk]);
        end
        if (PRED60_23_buffer[clk] != PRED60_23_buffer[!clk]) begin
          $fwrite(f, "Register (60,23) Value: %h\n", PRED60_23_buffer[clk]);
        end
        if (PRED60_24_buffer[clk] != PRED60_24_buffer[!clk]) begin
          $fwrite(f, "Register (60,24) Value: %h\n", PRED60_24_buffer[clk]);
        end
        if (PRED60_25_buffer[clk] != PRED60_25_buffer[!clk]) begin
          $fwrite(f, "Register (60,25) Value: %h\n", PRED60_25_buffer[clk]);
        end
        if (PRED60_26_buffer[clk] != PRED60_26_buffer[!clk]) begin
          $fwrite(f, "Register (60,26) Value: %h\n", PRED60_26_buffer[clk]);
        end
        if (PRED60_27_buffer[clk] != PRED60_27_buffer[!clk]) begin
          $fwrite(f, "Register (60,27) Value: %h\n", PRED60_27_buffer[clk]);
        end
        if (PRED60_28_buffer[clk] != PRED60_28_buffer[!clk]) begin
          $fwrite(f, "Register (60,28) Value: %h\n", PRED60_28_buffer[clk]);
        end
        if (PRED60_29_buffer[clk] != PRED60_29_buffer[!clk]) begin
          $fwrite(f, "Register (60,29) Value: %h\n", PRED60_29_buffer[clk]);
        end
        if (PRED60_30_buffer[clk] != PRED60_30_buffer[!clk]) begin
          $fwrite(f, "Register (60,30) Value: %h\n", PRED60_30_buffer[clk]);
        end
        if (PRED60_31_buffer[clk] != PRED60_31_buffer[!clk]) begin
          $fwrite(f, "Register (60,31) Value: %h\n", PRED60_31_buffer[clk]);
        end
        if (PRED61_0_buffer[clk] != PRED61_0_buffer[!clk]) begin
          $fwrite(f, "Register (61,0) Value: %h\n", PRED61_0_buffer[clk]);
        end
        if (PRED61_1_buffer[clk] != PRED61_1_buffer[!clk]) begin
          $fwrite(f, "Register (61,1) Value: %h\n", PRED61_1_buffer[clk]);
        end
        if (PRED61_2_buffer[clk] != PRED61_2_buffer[!clk]) begin
          $fwrite(f, "Register (61,2) Value: %h\n", PRED61_2_buffer[clk]);
        end
        if (PRED61_3_buffer[clk] != PRED61_3_buffer[!clk]) begin
          $fwrite(f, "Register (61,3) Value: %h\n", PRED61_3_buffer[clk]);
        end
        if (PRED61_4_buffer[clk] != PRED61_4_buffer[!clk]) begin
          $fwrite(f, "Register (61,4) Value: %h\n", PRED61_4_buffer[clk]);
        end
        if (PRED61_5_buffer[clk] != PRED61_5_buffer[!clk]) begin
          $fwrite(f, "Register (61,5) Value: %h\n", PRED61_5_buffer[clk]);
        end
        if (PRED61_6_buffer[clk] != PRED61_6_buffer[!clk]) begin
          $fwrite(f, "Register (61,6) Value: %h\n", PRED61_6_buffer[clk]);
        end
        if (PRED61_7_buffer[clk] != PRED61_7_buffer[!clk]) begin
          $fwrite(f, "Register (61,7) Value: %h\n", PRED61_7_buffer[clk]);
        end
        if (PRED61_8_buffer[clk] != PRED61_8_buffer[!clk]) begin
          $fwrite(f, "Register (61,8) Value: %h\n", PRED61_8_buffer[clk]);
        end
        if (PRED61_9_buffer[clk] != PRED61_9_buffer[!clk]) begin
          $fwrite(f, "Register (61,9) Value: %h\n", PRED61_9_buffer[clk]);
        end
        if (PRED61_10_buffer[clk] != PRED61_10_buffer[!clk]) begin
          $fwrite(f, "Register (61,10) Value: %h\n", PRED61_10_buffer[clk]);
        end
        if (PRED61_11_buffer[clk] != PRED61_11_buffer[!clk]) begin
          $fwrite(f, "Register (61,11) Value: %h\n", PRED61_11_buffer[clk]);
        end
        if (PRED61_12_buffer[clk] != PRED61_12_buffer[!clk]) begin
          $fwrite(f, "Register (61,12) Value: %h\n", PRED61_12_buffer[clk]);
        end
        if (PRED61_13_buffer[clk] != PRED61_13_buffer[!clk]) begin
          $fwrite(f, "Register (61,13) Value: %h\n", PRED61_13_buffer[clk]);
        end
        if (PRED61_14_buffer[clk] != PRED61_14_buffer[!clk]) begin
          $fwrite(f, "Register (61,14) Value: %h\n", PRED61_14_buffer[clk]);
        end
        if (PRED61_15_buffer[clk] != PRED61_15_buffer[!clk]) begin
          $fwrite(f, "Register (61,15) Value: %h\n", PRED61_15_buffer[clk]);
        end
        if (PRED61_16_buffer[clk] != PRED61_16_buffer[!clk]) begin
          $fwrite(f, "Register (61,16) Value: %h\n", PRED61_16_buffer[clk]);
        end
        if (PRED61_17_buffer[clk] != PRED61_17_buffer[!clk]) begin
          $fwrite(f, "Register (61,17) Value: %h\n", PRED61_17_buffer[clk]);
        end
        if (PRED61_18_buffer[clk] != PRED61_18_buffer[!clk]) begin
          $fwrite(f, "Register (61,18) Value: %h\n", PRED61_18_buffer[clk]);
        end
        if (PRED61_19_buffer[clk] != PRED61_19_buffer[!clk]) begin
          $fwrite(f, "Register (61,19) Value: %h\n", PRED61_19_buffer[clk]);
        end
        if (PRED61_20_buffer[clk] != PRED61_20_buffer[!clk]) begin
          $fwrite(f, "Register (61,20) Value: %h\n", PRED61_20_buffer[clk]);
        end
        if (PRED61_21_buffer[clk] != PRED61_21_buffer[!clk]) begin
          $fwrite(f, "Register (61,21) Value: %h\n", PRED61_21_buffer[clk]);
        end
        if (PRED61_22_buffer[clk] != PRED61_22_buffer[!clk]) begin
          $fwrite(f, "Register (61,22) Value: %h\n", PRED61_22_buffer[clk]);
        end
        if (PRED61_23_buffer[clk] != PRED61_23_buffer[!clk]) begin
          $fwrite(f, "Register (61,23) Value: %h\n", PRED61_23_buffer[clk]);
        end
        if (PRED61_24_buffer[clk] != PRED61_24_buffer[!clk]) begin
          $fwrite(f, "Register (61,24) Value: %h\n", PRED61_24_buffer[clk]);
        end
        if (PRED61_25_buffer[clk] != PRED61_25_buffer[!clk]) begin
          $fwrite(f, "Register (61,25) Value: %h\n", PRED61_25_buffer[clk]);
        end
        if (PRED61_26_buffer[clk] != PRED61_26_buffer[!clk]) begin
          $fwrite(f, "Register (61,26) Value: %h\n", PRED61_26_buffer[clk]);
        end
        if (PRED61_27_buffer[clk] != PRED61_27_buffer[!clk]) begin
          $fwrite(f, "Register (61,27) Value: %h\n", PRED61_27_buffer[clk]);
        end
        if (PRED61_28_buffer[clk] != PRED61_28_buffer[!clk]) begin
          $fwrite(f, "Register (61,28) Value: %h\n", PRED61_28_buffer[clk]);
        end
        if (PRED61_29_buffer[clk] != PRED61_29_buffer[!clk]) begin
          $fwrite(f, "Register (61,29) Value: %h\n", PRED61_29_buffer[clk]);
        end
        if (PRED61_30_buffer[clk] != PRED61_30_buffer[!clk]) begin
          $fwrite(f, "Register (61,30) Value: %h\n", PRED61_30_buffer[clk]);
        end
        if (PRED61_31_buffer[clk] != PRED61_31_buffer[!clk]) begin
          $fwrite(f, "Register (61,31) Value: %h\n", PRED61_31_buffer[clk]);
        end
        if (PRED62_0_buffer[clk] != PRED62_0_buffer[!clk]) begin
          $fwrite(f, "Register (62,0) Value: %h\n", PRED62_0_buffer[clk]);
        end
        if (PRED62_1_buffer[clk] != PRED62_1_buffer[!clk]) begin
          $fwrite(f, "Register (62,1) Value: %h\n", PRED62_1_buffer[clk]);
        end
        if (PRED62_2_buffer[clk] != PRED62_2_buffer[!clk]) begin
          $fwrite(f, "Register (62,2) Value: %h\n", PRED62_2_buffer[clk]);
        end
        if (PRED62_3_buffer[clk] != PRED62_3_buffer[!clk]) begin
          $fwrite(f, "Register (62,3) Value: %h\n", PRED62_3_buffer[clk]);
        end
        if (PRED62_4_buffer[clk] != PRED62_4_buffer[!clk]) begin
          $fwrite(f, "Register (62,4) Value: %h\n", PRED62_4_buffer[clk]);
        end
        if (PRED62_5_buffer[clk] != PRED62_5_buffer[!clk]) begin
          $fwrite(f, "Register (62,5) Value: %h\n", PRED62_5_buffer[clk]);
        end
        if (PRED62_6_buffer[clk] != PRED62_6_buffer[!clk]) begin
          $fwrite(f, "Register (62,6) Value: %h\n", PRED62_6_buffer[clk]);
        end
        if (PRED62_7_buffer[clk] != PRED62_7_buffer[!clk]) begin
          $fwrite(f, "Register (62,7) Value: %h\n", PRED62_7_buffer[clk]);
        end
        if (PRED62_8_buffer[clk] != PRED62_8_buffer[!clk]) begin
          $fwrite(f, "Register (62,8) Value: %h\n", PRED62_8_buffer[clk]);
        end
        if (PRED62_9_buffer[clk] != PRED62_9_buffer[!clk]) begin
          $fwrite(f, "Register (62,9) Value: %h\n", PRED62_9_buffer[clk]);
        end
        if (PRED62_10_buffer[clk] != PRED62_10_buffer[!clk]) begin
          $fwrite(f, "Register (62,10) Value: %h\n", PRED62_10_buffer[clk]);
        end
        if (PRED62_11_buffer[clk] != PRED62_11_buffer[!clk]) begin
          $fwrite(f, "Register (62,11) Value: %h\n", PRED62_11_buffer[clk]);
        end
        if (PRED62_12_buffer[clk] != PRED62_12_buffer[!clk]) begin
          $fwrite(f, "Register (62,12) Value: %h\n", PRED62_12_buffer[clk]);
        end
        if (PRED62_13_buffer[clk] != PRED62_13_buffer[!clk]) begin
          $fwrite(f, "Register (62,13) Value: %h\n", PRED62_13_buffer[clk]);
        end
        if (PRED62_14_buffer[clk] != PRED62_14_buffer[!clk]) begin
          $fwrite(f, "Register (62,14) Value: %h\n", PRED62_14_buffer[clk]);
        end
        if (PRED62_15_buffer[clk] != PRED62_15_buffer[!clk]) begin
          $fwrite(f, "Register (62,15) Value: %h\n", PRED62_15_buffer[clk]);
        end
        if (PRED62_16_buffer[clk] != PRED62_16_buffer[!clk]) begin
          $fwrite(f, "Register (62,16) Value: %h\n", PRED62_16_buffer[clk]);
        end
        if (PRED62_17_buffer[clk] != PRED62_17_buffer[!clk]) begin
          $fwrite(f, "Register (62,17) Value: %h\n", PRED62_17_buffer[clk]);
        end
        if (PRED62_18_buffer[clk] != PRED62_18_buffer[!clk]) begin
          $fwrite(f, "Register (62,18) Value: %h\n", PRED62_18_buffer[clk]);
        end
        if (PRED62_19_buffer[clk] != PRED62_19_buffer[!clk]) begin
          $fwrite(f, "Register (62,19) Value: %h\n", PRED62_19_buffer[clk]);
        end
        if (PRED62_20_buffer[clk] != PRED62_20_buffer[!clk]) begin
          $fwrite(f, "Register (62,20) Value: %h\n", PRED62_20_buffer[clk]);
        end
        if (PRED62_21_buffer[clk] != PRED62_21_buffer[!clk]) begin
          $fwrite(f, "Register (62,21) Value: %h\n", PRED62_21_buffer[clk]);
        end
        if (PRED62_22_buffer[clk] != PRED62_22_buffer[!clk]) begin
          $fwrite(f, "Register (62,22) Value: %h\n", PRED62_22_buffer[clk]);
        end
        if (PRED62_23_buffer[clk] != PRED62_23_buffer[!clk]) begin
          $fwrite(f, "Register (62,23) Value: %h\n", PRED62_23_buffer[clk]);
        end
        if (PRED62_24_buffer[clk] != PRED62_24_buffer[!clk]) begin
          $fwrite(f, "Register (62,24) Value: %h\n", PRED62_24_buffer[clk]);
        end
        if (PRED62_25_buffer[clk] != PRED62_25_buffer[!clk]) begin
          $fwrite(f, "Register (62,25) Value: %h\n", PRED62_25_buffer[clk]);
        end
        if (PRED62_26_buffer[clk] != PRED62_26_buffer[!clk]) begin
          $fwrite(f, "Register (62,26) Value: %h\n", PRED62_26_buffer[clk]);
        end
        if (PRED62_27_buffer[clk] != PRED62_27_buffer[!clk]) begin
          $fwrite(f, "Register (62,27) Value: %h\n", PRED62_27_buffer[clk]);
        end
        if (PRED62_28_buffer[clk] != PRED62_28_buffer[!clk]) begin
          $fwrite(f, "Register (62,28) Value: %h\n", PRED62_28_buffer[clk]);
        end
        if (PRED62_29_buffer[clk] != PRED62_29_buffer[!clk]) begin
          $fwrite(f, "Register (62,29) Value: %h\n", PRED62_29_buffer[clk]);
        end
        if (PRED62_30_buffer[clk] != PRED62_30_buffer[!clk]) begin
          $fwrite(f, "Register (62,30) Value: %h\n", PRED62_30_buffer[clk]);
        end
        if (PRED62_31_buffer[clk] != PRED62_31_buffer[!clk]) begin
          $fwrite(f, "Register (62,31) Value: %h\n", PRED62_31_buffer[clk]);
        end
        if (PRED63_0_buffer[clk] != PRED63_0_buffer[!clk]) begin
          $fwrite(f, "Register (63,0) Value: %h\n", PRED63_0_buffer[clk]);
        end
        if (PRED63_1_buffer[clk] != PRED63_1_buffer[!clk]) begin
          $fwrite(f, "Register (63,1) Value: %h\n", PRED63_1_buffer[clk]);
        end
        if (PRED63_2_buffer[clk] != PRED63_2_buffer[!clk]) begin
          $fwrite(f, "Register (63,2) Value: %h\n", PRED63_2_buffer[clk]);
        end
        if (PRED63_3_buffer[clk] != PRED63_3_buffer[!clk]) begin
          $fwrite(f, "Register (63,3) Value: %h\n", PRED63_3_buffer[clk]);
        end
        if (PRED63_4_buffer[clk] != PRED63_4_buffer[!clk]) begin
          $fwrite(f, "Register (63,4) Value: %h\n", PRED63_4_buffer[clk]);
        end
        if (PRED63_5_buffer[clk] != PRED63_5_buffer[!clk]) begin
          $fwrite(f, "Register (63,5) Value: %h\n", PRED63_5_buffer[clk]);
        end
        if (PRED63_6_buffer[clk] != PRED63_6_buffer[!clk]) begin
          $fwrite(f, "Register (63,6) Value: %h\n", PRED63_6_buffer[clk]);
        end
        if (PRED63_7_buffer[clk] != PRED63_7_buffer[!clk]) begin
          $fwrite(f, "Register (63,7) Value: %h\n", PRED63_7_buffer[clk]);
        end
        if (PRED63_8_buffer[clk] != PRED63_8_buffer[!clk]) begin
          $fwrite(f, "Register (63,8) Value: %h\n", PRED63_8_buffer[clk]);
        end
        if (PRED63_9_buffer[clk] != PRED63_9_buffer[!clk]) begin
          $fwrite(f, "Register (63,9) Value: %h\n", PRED63_9_buffer[clk]);
        end
        if (PRED63_10_buffer[clk] != PRED63_10_buffer[!clk]) begin
          $fwrite(f, "Register (63,10) Value: %h\n", PRED63_10_buffer[clk]);
        end
        if (PRED63_11_buffer[clk] != PRED63_11_buffer[!clk]) begin
          $fwrite(f, "Register (63,11) Value: %h\n", PRED63_11_buffer[clk]);
        end
        if (PRED63_12_buffer[clk] != PRED63_12_buffer[!clk]) begin
          $fwrite(f, "Register (63,12) Value: %h\n", PRED63_12_buffer[clk]);
        end
        if (PRED63_13_buffer[clk] != PRED63_13_buffer[!clk]) begin
          $fwrite(f, "Register (63,13) Value: %h\n", PRED63_13_buffer[clk]);
        end
        if (PRED63_14_buffer[clk] != PRED63_14_buffer[!clk]) begin
          $fwrite(f, "Register (63,14) Value: %h\n", PRED63_14_buffer[clk]);
        end
        if (PRED63_15_buffer[clk] != PRED63_15_buffer[!clk]) begin
          $fwrite(f, "Register (63,15) Value: %h\n", PRED63_15_buffer[clk]);
        end
        if (PRED63_16_buffer[clk] != PRED63_16_buffer[!clk]) begin
          $fwrite(f, "Register (63,16) Value: %h\n", PRED63_16_buffer[clk]);
        end
        if (PRED63_17_buffer[clk] != PRED63_17_buffer[!clk]) begin
          $fwrite(f, "Register (63,17) Value: %h\n", PRED63_17_buffer[clk]);
        end
        if (PRED63_18_buffer[clk] != PRED63_18_buffer[!clk]) begin
          $fwrite(f, "Register (63,18) Value: %h\n", PRED63_18_buffer[clk]);
        end
        if (PRED63_19_buffer[clk] != PRED63_19_buffer[!clk]) begin
          $fwrite(f, "Register (63,19) Value: %h\n", PRED63_19_buffer[clk]);
        end
        if (PRED63_20_buffer[clk] != PRED63_20_buffer[!clk]) begin
          $fwrite(f, "Register (63,20) Value: %h\n", PRED63_20_buffer[clk]);
        end
        if (PRED63_21_buffer[clk] != PRED63_21_buffer[!clk]) begin
          $fwrite(f, "Register (63,21) Value: %h\n", PRED63_21_buffer[clk]);
        end
        if (PRED63_22_buffer[clk] != PRED63_22_buffer[!clk]) begin
          $fwrite(f, "Register (63,22) Value: %h\n", PRED63_22_buffer[clk]);
        end
        if (PRED63_23_buffer[clk] != PRED63_23_buffer[!clk]) begin
          $fwrite(f, "Register (63,23) Value: %h\n", PRED63_23_buffer[clk]);
        end
        if (PRED63_24_buffer[clk] != PRED63_24_buffer[!clk]) begin
          $fwrite(f, "Register (63,24) Value: %h\n", PRED63_24_buffer[clk]);
        end
        if (PRED63_25_buffer[clk] != PRED63_25_buffer[!clk]) begin
          $fwrite(f, "Register (63,25) Value: %h\n", PRED63_25_buffer[clk]);
        end
        if (PRED63_26_buffer[clk] != PRED63_26_buffer[!clk]) begin
          $fwrite(f, "Register (63,26) Value: %h\n", PRED63_26_buffer[clk]);
        end
        if (PRED63_27_buffer[clk] != PRED63_27_buffer[!clk]) begin
          $fwrite(f, "Register (63,27) Value: %h\n", PRED63_27_buffer[clk]);
        end
        if (PRED63_28_buffer[clk] != PRED63_28_buffer[!clk]) begin
          $fwrite(f, "Register (63,28) Value: %h\n", PRED63_28_buffer[clk]);
        end
        if (PRED63_29_buffer[clk] != PRED63_29_buffer[!clk]) begin
          $fwrite(f, "Register (63,29) Value: %h\n", PRED63_29_buffer[clk]);
        end
        if (PRED63_30_buffer[clk] != PRED63_30_buffer[!clk]) begin
          $fwrite(f, "Register (63,30) Value: %h\n", PRED63_30_buffer[clk]);
        end
        if (PRED63_31_buffer[clk] != PRED63_31_buffer[!clk]) begin
          $fwrite(f, "Register (63,31) Value: %h\n", PRED63_31_buffer[clk]);
        end

        $fwrite(f, " \n=====================================================\n\n\n\n\n");
      end
    end
    $fclose(f);
  end 

endmodule









