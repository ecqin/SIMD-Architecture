//===================================================================
// Filename: harmonica_tracker.sv
// Author: Eric Qin
// Purpose: Verification Module (test debugger)
//===================================================================


// Under Development
// TODO List
// 1) MACRO to get essential values in a readable form (non-synthesizable) // TODO
// 2) Print out of the register files based on thre warp and thread ID to read
// 3) Also serves as a checker and print out potential failed cases and timestamp
// 4) Look into tasks and interfaces
// 5) Make it generic to the point that timing changes doesnt affect the output as much
// FIXME -> code structure not efficient, too lengthy


`include "harmonica_cfg.sv" 

module harmonica_tracker(
  input logic clk,
  // FIXME --> very wordy, not efficient
  // Interfaces? tasks? structs? need to look into this in the future
/*
  generate
    genvar GPR_index;
    for (GPR_index=0; GPR_index<NUM_TOTAL_THREADS; GPR_index=GPR_index+1) begin
      input logic [63:0] .NAME("GPR" + GPR_index)  [0:31];
    end
  endgenerate
*/
  input logic [63:0] GRF0 [0:31],
  input logic [63:0] GRF1 [0:31],
  input logic [63:0] GRF2 [0:31],
  input logic [63:0] GRF3 [0:31],
  input logic [63:0] GRF4 [0:31],
  input logic [63:0] GRF5 [0:31],
  input logic [63:0] GRF6 [0:31],
  input logic [63:0] GRF7 [0:31],
  input logic [63:0] GRF8 [0:31],
  input logic [63:0] GRF9 [0:31],
  input logic [63:0] GRF10 [0:31],
  input logic [63:0] GRF11 [0:31],
  input logic [63:0] GRF12 [0:31],
  input logic [63:0] GRF13 [0:31],
  input logic [63:0] GRF14 [0:31],
  input logic [63:0] GRF15 [0:31],
  input logic [63:0] GRF16 [0:31],
  input logic [63:0] GRF17 [0:31],
  input logic [63:0] GRF18 [0:31],
  input logic [63:0] GRF19 [0:31],
  input logic [63:0] GRF20 [0:31],
  input logic [63:0] GRF21 [0:31],
  input logic [63:0] GRF22 [0:31],
  input logic [63:0] GRF23 [0:31],
  input logic [63:0] GRF24 [0:31],
  input logic [63:0] GRF25 [0:31],
  input logic [63:0] GRF26 [0:31],
  input logic [63:0] GRF27 [0:31],
  input logic [63:0] GRF28 [0:31],
  input logic [63:0] GRF29 [0:31],
  input logic [63:0] GRF30 [0:31],
  input logic [63:0] GRF31 [0:31],
  input logic [63:0] GRF32 [0:31],
  input logic [63:0] GRF33 [0:31],
  input logic [63:0] GRF34 [0:31],
  input logic [63:0] GRF35 [0:31],
  input logic [63:0] GRF36 [0:31],
  input logic [63:0] GRF37 [0:31],
  input logic [63:0] GRF38 [0:31],
  input logic [63:0] GRF39 [0:31],
  input logic [63:0] GRF40 [0:31],
  input logic [63:0] GRF41 [0:31],
  input logic [63:0] GRF42 [0:31],
  input logic [63:0] GRF43 [0:31],
  input logic [63:0] GRF44 [0:31],
  input logic [63:0] GRF45 [0:31],
  input logic [63:0] GRF46 [0:31],
  input logic [63:0] GRF47 [0:31],
  input logic [63:0] GRF48 [0:31],
  input logic [63:0] GRF49 [0:31],
  input logic [63:0] GRF50 [0:31],
  input logic [63:0] GRF51 [0:31],
  input logic [63:0] GRF52 [0:31],
  input logic [63:0] GRF53 [0:31],
  input logic [63:0] GRF54 [0:31],
  input logic [63:0] GRF55 [0:31],
  input logic [63:0] GRF56 [0:31],
  input logic [63:0] GRF57 [0:31],
  input logic [63:0] GRF58 [0:31],
  input logic [63:0] GRF59 [0:31],
  input logic [63:0] GRF60 [0:31],
  input logic [63:0] GRF61 [0:31],
  input logic [63:0] GRF62 [0:31],
  input logic [63:0] GRF63 [0:31]
);

  integer f, i;
  // Initialize 2-entry buffers for comparison....

  // All register entry in all register files, code bloat. FIXME please, must be a better way, genvar???? 
  // 64 * 32 lol........
  logic [63:0] GRF0_0_buffer [0:1];
  logic [63:0] GRF0_1_buffer [0:1];
  logic [63:0] GRF0_2_buffer [0:1];
  logic [63:0] GRF0_3_buffer [0:1];
  logic [63:0] GRF0_4_buffer [0:1];
  logic [63:0] GRF0_5_buffer [0:1];
  logic [63:0] GRF0_6_buffer [0:1];
  logic [63:0] GRF0_7_buffer [0:1];
  logic [63:0] GRF0_8_buffer [0:1];
  logic [63:0] GRF0_9_buffer [0:1];
  logic [63:0] GRF0_10_buffer [0:1];
  logic [63:0] GRF0_11_buffer [0:1];
  logic [63:0] GRF0_12_buffer [0:1];
  logic [63:0] GRF0_13_buffer [0:1];
  logic [63:0] GRF0_14_buffer [0:1];
  logic [63:0] GRF0_15_buffer [0:1];
  logic [63:0] GRF0_16_buffer [0:1];
  logic [63:0] GRF0_17_buffer [0:1];
  logic [63:0] GRF0_18_buffer [0:1];
  logic [63:0] GRF0_19_buffer [0:1];
  logic [63:0] GRF0_20_buffer [0:1];
  logic [63:0] GRF0_21_buffer [0:1];
  logic [63:0] GRF0_22_buffer [0:1];
  logic [63:0] GRF0_23_buffer [0:1];
  logic [63:0] GRF0_24_buffer [0:1];
  logic [63:0] GRF0_25_buffer [0:1];
  logic [63:0] GRF0_26_buffer [0:1];
  logic [63:0] GRF0_27_buffer [0:1];
  logic [63:0] GRF0_28_buffer [0:1];
  logic [63:0] GRF0_29_buffer [0:1];
  logic [63:0] GRF0_30_buffer [0:1];
  logic [63:0] GRF0_31_buffer [0:1];
  logic [63:0] GRF1_0_buffer [0:1];
  logic [63:0] GRF1_1_buffer [0:1];
  logic [63:0] GRF1_2_buffer [0:1];
  logic [63:0] GRF1_3_buffer [0:1];
  logic [63:0] GRF1_4_buffer [0:1];
  logic [63:0] GRF1_5_buffer [0:1];
  logic [63:0] GRF1_6_buffer [0:1];
  logic [63:0] GRF1_7_buffer [0:1];
  logic [63:0] GRF1_8_buffer [0:1];
  logic [63:0] GRF1_9_buffer [0:1];
  logic [63:0] GRF1_10_buffer [0:1];
  logic [63:0] GRF1_11_buffer [0:1];
  logic [63:0] GRF1_12_buffer [0:1];
  logic [63:0] GRF1_13_buffer [0:1];
  logic [63:0] GRF1_14_buffer [0:1];
  logic [63:0] GRF1_15_buffer [0:1];
  logic [63:0] GRF1_16_buffer [0:1];
  logic [63:0] GRF1_17_buffer [0:1];
  logic [63:0] GRF1_18_buffer [0:1];
  logic [63:0] GRF1_19_buffer [0:1];
  logic [63:0] GRF1_20_buffer [0:1];
  logic [63:0] GRF1_21_buffer [0:1];
  logic [63:0] GRF1_22_buffer [0:1];
  logic [63:0] GRF1_23_buffer [0:1];
  logic [63:0] GRF1_24_buffer [0:1];
  logic [63:0] GRF1_25_buffer [0:1];
  logic [63:0] GRF1_26_buffer [0:1];
  logic [63:0] GRF1_27_buffer [0:1];
  logic [63:0] GRF1_28_buffer [0:1];
  logic [63:0] GRF1_29_buffer [0:1];
  logic [63:0] GRF1_30_buffer [0:1];
  logic [63:0] GRF1_31_buffer [0:1];
  logic [63:0] GRF2_0_buffer [0:1];
  logic [63:0] GRF2_1_buffer [0:1];
  logic [63:0] GRF2_2_buffer [0:1];
  logic [63:0] GRF2_3_buffer [0:1];
  logic [63:0] GRF2_4_buffer [0:1];
  logic [63:0] GRF2_5_buffer [0:1];
  logic [63:0] GRF2_6_buffer [0:1];
  logic [63:0] GRF2_7_buffer [0:1];
  logic [63:0] GRF2_8_buffer [0:1];
  logic [63:0] GRF2_9_buffer [0:1];
  logic [63:0] GRF2_10_buffer [0:1];
  logic [63:0] GRF2_11_buffer [0:1];
  logic [63:0] GRF2_12_buffer [0:1];
  logic [63:0] GRF2_13_buffer [0:1];
  logic [63:0] GRF2_14_buffer [0:1];
  logic [63:0] GRF2_15_buffer [0:1];
  logic [63:0] GRF2_16_buffer [0:1];
  logic [63:0] GRF2_17_buffer [0:1];
  logic [63:0] GRF2_18_buffer [0:1];
  logic [63:0] GRF2_19_buffer [0:1];
  logic [63:0] GRF2_20_buffer [0:1];
  logic [63:0] GRF2_21_buffer [0:1];
  logic [63:0] GRF2_22_buffer [0:1];
  logic [63:0] GRF2_23_buffer [0:1];
  logic [63:0] GRF2_24_buffer [0:1];
  logic [63:0] GRF2_25_buffer [0:1];
  logic [63:0] GRF2_26_buffer [0:1];
  logic [63:0] GRF2_27_buffer [0:1];
  logic [63:0] GRF2_28_buffer [0:1];
  logic [63:0] GRF2_29_buffer [0:1];
  logic [63:0] GRF2_30_buffer [0:1];
  logic [63:0] GRF2_31_buffer [0:1];
  logic [63:0] GRF3_0_buffer [0:1];
  logic [63:0] GRF3_1_buffer [0:1];
  logic [63:0] GRF3_2_buffer [0:1];
  logic [63:0] GRF3_3_buffer [0:1];
  logic [63:0] GRF3_4_buffer [0:1];
  logic [63:0] GRF3_5_buffer [0:1];
  logic [63:0] GRF3_6_buffer [0:1];
  logic [63:0] GRF3_7_buffer [0:1];
  logic [63:0] GRF3_8_buffer [0:1];
  logic [63:0] GRF3_9_buffer [0:1];
  logic [63:0] GRF3_10_buffer [0:1];
  logic [63:0] GRF3_11_buffer [0:1];
  logic [63:0] GRF3_12_buffer [0:1];
  logic [63:0] GRF3_13_buffer [0:1];
  logic [63:0] GRF3_14_buffer [0:1];
  logic [63:0] GRF3_15_buffer [0:1];
  logic [63:0] GRF3_16_buffer [0:1];
  logic [63:0] GRF3_17_buffer [0:1];
  logic [63:0] GRF3_18_buffer [0:1];
  logic [63:0] GRF3_19_buffer [0:1];
  logic [63:0] GRF3_20_buffer [0:1];
  logic [63:0] GRF3_21_buffer [0:1];
  logic [63:0] GRF3_22_buffer [0:1];
  logic [63:0] GRF3_23_buffer [0:1];
  logic [63:0] GRF3_24_buffer [0:1];
  logic [63:0] GRF3_25_buffer [0:1];
  logic [63:0] GRF3_26_buffer [0:1];
  logic [63:0] GRF3_27_buffer [0:1];
  logic [63:0] GRF3_28_buffer [0:1];
  logic [63:0] GRF3_29_buffer [0:1];
  logic [63:0] GRF3_30_buffer [0:1];
  logic [63:0] GRF3_31_buffer [0:1];
  logic [63:0] GRF4_0_buffer [0:1];
  logic [63:0] GRF4_1_buffer [0:1];
  logic [63:0] GRF4_2_buffer [0:1];
  logic [63:0] GRF4_3_buffer [0:1];
  logic [63:0] GRF4_4_buffer [0:1];
  logic [63:0] GRF4_5_buffer [0:1];
  logic [63:0] GRF4_6_buffer [0:1];
  logic [63:0] GRF4_7_buffer [0:1];
  logic [63:0] GRF4_8_buffer [0:1];
  logic [63:0] GRF4_9_buffer [0:1];
  logic [63:0] GRF4_10_buffer [0:1];
  logic [63:0] GRF4_11_buffer [0:1];
  logic [63:0] GRF4_12_buffer [0:1];
  logic [63:0] GRF4_13_buffer [0:1];
  logic [63:0] GRF4_14_buffer [0:1];
  logic [63:0] GRF4_15_buffer [0:1];
  logic [63:0] GRF4_16_buffer [0:1];
  logic [63:0] GRF4_17_buffer [0:1];
  logic [63:0] GRF4_18_buffer [0:1];
  logic [63:0] GRF4_19_buffer [0:1];
  logic [63:0] GRF4_20_buffer [0:1];
  logic [63:0] GRF4_21_buffer [0:1];
  logic [63:0] GRF4_22_buffer [0:1];
  logic [63:0] GRF4_23_buffer [0:1];
  logic [63:0] GRF4_24_buffer [0:1];
  logic [63:0] GRF4_25_buffer [0:1];
  logic [63:0] GRF4_26_buffer [0:1];
  logic [63:0] GRF4_27_buffer [0:1];
  logic [63:0] GRF4_28_buffer [0:1];
  logic [63:0] GRF4_29_buffer [0:1];
  logic [63:0] GRF4_30_buffer [0:1];
  logic [63:0] GRF4_31_buffer [0:1];
  logic [63:0] GRF5_0_buffer [0:1];
  logic [63:0] GRF5_1_buffer [0:1];
  logic [63:0] GRF5_2_buffer [0:1];
  logic [63:0] GRF5_3_buffer [0:1];
  logic [63:0] GRF5_4_buffer [0:1];
  logic [63:0] GRF5_5_buffer [0:1];
  logic [63:0] GRF5_6_buffer [0:1];
  logic [63:0] GRF5_7_buffer [0:1];
  logic [63:0] GRF5_8_buffer [0:1];
  logic [63:0] GRF5_9_buffer [0:1];
  logic [63:0] GRF5_10_buffer [0:1];
  logic [63:0] GRF5_11_buffer [0:1];
  logic [63:0] GRF5_12_buffer [0:1];
  logic [63:0] GRF5_13_buffer [0:1];
  logic [63:0] GRF5_14_buffer [0:1];
  logic [63:0] GRF5_15_buffer [0:1];
  logic [63:0] GRF5_16_buffer [0:1];
  logic [63:0] GRF5_17_buffer [0:1];
  logic [63:0] GRF5_18_buffer [0:1];
  logic [63:0] GRF5_19_buffer [0:1];
  logic [63:0] GRF5_20_buffer [0:1];
  logic [63:0] GRF5_21_buffer [0:1];
  logic [63:0] GRF5_22_buffer [0:1];
  logic [63:0] GRF5_23_buffer [0:1];
  logic [63:0] GRF5_24_buffer [0:1];
  logic [63:0] GRF5_25_buffer [0:1];
  logic [63:0] GRF5_26_buffer [0:1];
  logic [63:0] GRF5_27_buffer [0:1];
  logic [63:0] GRF5_28_buffer [0:1];
  logic [63:0] GRF5_29_buffer [0:1];
  logic [63:0] GRF5_30_buffer [0:1];
  logic [63:0] GRF5_31_buffer [0:1];
  logic [63:0] GRF6_0_buffer [0:1];
  logic [63:0] GRF6_1_buffer [0:1];
  logic [63:0] GRF6_2_buffer [0:1];
  logic [63:0] GRF6_3_buffer [0:1];
  logic [63:0] GRF6_4_buffer [0:1];
  logic [63:0] GRF6_5_buffer [0:1];
  logic [63:0] GRF6_6_buffer [0:1];
  logic [63:0] GRF6_7_buffer [0:1];
  logic [63:0] GRF6_8_buffer [0:1];
  logic [63:0] GRF6_9_buffer [0:1];
  logic [63:0] GRF6_10_buffer [0:1];
  logic [63:0] GRF6_11_buffer [0:1];
  logic [63:0] GRF6_12_buffer [0:1];
  logic [63:0] GRF6_13_buffer [0:1];
  logic [63:0] GRF6_14_buffer [0:1];
  logic [63:0] GRF6_15_buffer [0:1];
  logic [63:0] GRF6_16_buffer [0:1];
  logic [63:0] GRF6_17_buffer [0:1];
  logic [63:0] GRF6_18_buffer [0:1];
  logic [63:0] GRF6_19_buffer [0:1];
  logic [63:0] GRF6_20_buffer [0:1];
  logic [63:0] GRF6_21_buffer [0:1];
  logic [63:0] GRF6_22_buffer [0:1];
  logic [63:0] GRF6_23_buffer [0:1];
  logic [63:0] GRF6_24_buffer [0:1];
  logic [63:0] GRF6_25_buffer [0:1];
  logic [63:0] GRF6_26_buffer [0:1];
  logic [63:0] GRF6_27_buffer [0:1];
  logic [63:0] GRF6_28_buffer [0:1];
  logic [63:0] GRF6_29_buffer [0:1];
  logic [63:0] GRF6_30_buffer [0:1];
  logic [63:0] GRF6_31_buffer [0:1];
  logic [63:0] GRF7_0_buffer [0:1];
  logic [63:0] GRF7_1_buffer [0:1];
  logic [63:0] GRF7_2_buffer [0:1];
  logic [63:0] GRF7_3_buffer [0:1];
  logic [63:0] GRF7_4_buffer [0:1];
  logic [63:0] GRF7_5_buffer [0:1];
  logic [63:0] GRF7_6_buffer [0:1];
  logic [63:0] GRF7_7_buffer [0:1];
  logic [63:0] GRF7_8_buffer [0:1];
  logic [63:0] GRF7_9_buffer [0:1];
  logic [63:0] GRF7_10_buffer [0:1];
  logic [63:0] GRF7_11_buffer [0:1];
  logic [63:0] GRF7_12_buffer [0:1];
  logic [63:0] GRF7_13_buffer [0:1];
  logic [63:0] GRF7_14_buffer [0:1];
  logic [63:0] GRF7_15_buffer [0:1];
  logic [63:0] GRF7_16_buffer [0:1];
  logic [63:0] GRF7_17_buffer [0:1];
  logic [63:0] GRF7_18_buffer [0:1];
  logic [63:0] GRF7_19_buffer [0:1];
  logic [63:0] GRF7_20_buffer [0:1];
  logic [63:0] GRF7_21_buffer [0:1];
  logic [63:0] GRF7_22_buffer [0:1];
  logic [63:0] GRF7_23_buffer [0:1];
  logic [63:0] GRF7_24_buffer [0:1];
  logic [63:0] GRF7_25_buffer [0:1];
  logic [63:0] GRF7_26_buffer [0:1];
  logic [63:0] GRF7_27_buffer [0:1];
  logic [63:0] GRF7_28_buffer [0:1];
  logic [63:0] GRF7_29_buffer [0:1];
  logic [63:0] GRF7_30_buffer [0:1];
  logic [63:0] GRF7_31_buffer [0:1];
  logic [63:0] GRF8_0_buffer [0:1];
  logic [63:0] GRF8_1_buffer [0:1];
  logic [63:0] GRF8_2_buffer [0:1];
  logic [63:0] GRF8_3_buffer [0:1];
  logic [63:0] GRF8_4_buffer [0:1];
  logic [63:0] GRF8_5_buffer [0:1];
  logic [63:0] GRF8_6_buffer [0:1];
  logic [63:0] GRF8_7_buffer [0:1];
  logic [63:0] GRF8_8_buffer [0:1];
  logic [63:0] GRF8_9_buffer [0:1];
  logic [63:0] GRF8_10_buffer [0:1];
  logic [63:0] GRF8_11_buffer [0:1];
  logic [63:0] GRF8_12_buffer [0:1];
  logic [63:0] GRF8_13_buffer [0:1];
  logic [63:0] GRF8_14_buffer [0:1];
  logic [63:0] GRF8_15_buffer [0:1];
  logic [63:0] GRF8_16_buffer [0:1];
  logic [63:0] GRF8_17_buffer [0:1];
  logic [63:0] GRF8_18_buffer [0:1];
  logic [63:0] GRF8_19_buffer [0:1];
  logic [63:0] GRF8_20_buffer [0:1];
  logic [63:0] GRF8_21_buffer [0:1];
  logic [63:0] GRF8_22_buffer [0:1];
  logic [63:0] GRF8_23_buffer [0:1];
  logic [63:0] GRF8_24_buffer [0:1];
  logic [63:0] GRF8_25_buffer [0:1];
  logic [63:0] GRF8_26_buffer [0:1];
  logic [63:0] GRF8_27_buffer [0:1];
  logic [63:0] GRF8_28_buffer [0:1];
  logic [63:0] GRF8_29_buffer [0:1];
  logic [63:0] GRF8_30_buffer [0:1];
  logic [63:0] GRF8_31_buffer [0:1];
  logic [63:0] GRF9_0_buffer [0:1];
  logic [63:0] GRF9_1_buffer [0:1];
  logic [63:0] GRF9_2_buffer [0:1];
  logic [63:0] GRF9_3_buffer [0:1];
  logic [63:0] GRF9_4_buffer [0:1];
  logic [63:0] GRF9_5_buffer [0:1];
  logic [63:0] GRF9_6_buffer [0:1];
  logic [63:0] GRF9_7_buffer [0:1];
  logic [63:0] GRF9_8_buffer [0:1];
  logic [63:0] GRF9_9_buffer [0:1];
  logic [63:0] GRF9_10_buffer [0:1];
  logic [63:0] GRF9_11_buffer [0:1];
  logic [63:0] GRF9_12_buffer [0:1];
  logic [63:0] GRF9_13_buffer [0:1];
  logic [63:0] GRF9_14_buffer [0:1];
  logic [63:0] GRF9_15_buffer [0:1];
  logic [63:0] GRF9_16_buffer [0:1];
  logic [63:0] GRF9_17_buffer [0:1];
  logic [63:0] GRF9_18_buffer [0:1];
  logic [63:0] GRF9_19_buffer [0:1];
  logic [63:0] GRF9_20_buffer [0:1];
  logic [63:0] GRF9_21_buffer [0:1];
  logic [63:0] GRF9_22_buffer [0:1];
  logic [63:0] GRF9_23_buffer [0:1];
  logic [63:0] GRF9_24_buffer [0:1];
  logic [63:0] GRF9_25_buffer [0:1];
  logic [63:0] GRF9_26_buffer [0:1];
  logic [63:0] GRF9_27_buffer [0:1];
  logic [63:0] GRF9_28_buffer [0:1];
  logic [63:0] GRF9_29_buffer [0:1];
  logic [63:0] GRF9_30_buffer [0:1];
  logic [63:0] GRF9_31_buffer [0:1];
  logic [63:0] GRF10_0_buffer [0:1];
  logic [63:0] GRF10_1_buffer [0:1];
  logic [63:0] GRF10_2_buffer [0:1];
  logic [63:0] GRF10_3_buffer [0:1];
  logic [63:0] GRF10_4_buffer [0:1];
  logic [63:0] GRF10_5_buffer [0:1];
  logic [63:0] GRF10_6_buffer [0:1];
  logic [63:0] GRF10_7_buffer [0:1];
  logic [63:0] GRF10_8_buffer [0:1];
  logic [63:0] GRF10_9_buffer [0:1];
  logic [63:0] GRF10_10_buffer [0:1];
  logic [63:0] GRF10_11_buffer [0:1];
  logic [63:0] GRF10_12_buffer [0:1];
  logic [63:0] GRF10_13_buffer [0:1];
  logic [63:0] GRF10_14_buffer [0:1];
  logic [63:0] GRF10_15_buffer [0:1];
  logic [63:0] GRF10_16_buffer [0:1];
  logic [63:0] GRF10_17_buffer [0:1];
  logic [63:0] GRF10_18_buffer [0:1];
  logic [63:0] GRF10_19_buffer [0:1];
  logic [63:0] GRF10_20_buffer [0:1];
  logic [63:0] GRF10_21_buffer [0:1];
  logic [63:0] GRF10_22_buffer [0:1];
  logic [63:0] GRF10_23_buffer [0:1];
  logic [63:0] GRF10_24_buffer [0:1];
  logic [63:0] GRF10_25_buffer [0:1];
  logic [63:0] GRF10_26_buffer [0:1];
  logic [63:0] GRF10_27_buffer [0:1];
  logic [63:0] GRF10_28_buffer [0:1];
  logic [63:0] GRF10_29_buffer [0:1];
  logic [63:0] GRF10_30_buffer [0:1];
  logic [63:0] GRF10_31_buffer [0:1];
  logic [63:0] GRF11_0_buffer [0:1];
  logic [63:0] GRF11_1_buffer [0:1];
  logic [63:0] GRF11_2_buffer [0:1];
  logic [63:0] GRF11_3_buffer [0:1];
  logic [63:0] GRF11_4_buffer [0:1];
  logic [63:0] GRF11_5_buffer [0:1];
  logic [63:0] GRF11_6_buffer [0:1];
  logic [63:0] GRF11_7_buffer [0:1];
  logic [63:0] GRF11_8_buffer [0:1];
  logic [63:0] GRF11_9_buffer [0:1];
  logic [63:0] GRF11_10_buffer [0:1];
  logic [63:0] GRF11_11_buffer [0:1];
  logic [63:0] GRF11_12_buffer [0:1];
  logic [63:0] GRF11_13_buffer [0:1];
  logic [63:0] GRF11_14_buffer [0:1];
  logic [63:0] GRF11_15_buffer [0:1];
  logic [63:0] GRF11_16_buffer [0:1];
  logic [63:0] GRF11_17_buffer [0:1];
  logic [63:0] GRF11_18_buffer [0:1];
  logic [63:0] GRF11_19_buffer [0:1];
  logic [63:0] GRF11_20_buffer [0:1];
  logic [63:0] GRF11_21_buffer [0:1];
  logic [63:0] GRF11_22_buffer [0:1];
  logic [63:0] GRF11_23_buffer [0:1];
  logic [63:0] GRF11_24_buffer [0:1];
  logic [63:0] GRF11_25_buffer [0:1];
  logic [63:0] GRF11_26_buffer [0:1];
  logic [63:0] GRF11_27_buffer [0:1];
  logic [63:0] GRF11_28_buffer [0:1];
  logic [63:0] GRF11_29_buffer [0:1];
  logic [63:0] GRF11_30_buffer [0:1];
  logic [63:0] GRF11_31_buffer [0:1];
  logic [63:0] GRF12_0_buffer [0:1];
  logic [63:0] GRF12_1_buffer [0:1];
  logic [63:0] GRF12_2_buffer [0:1];
  logic [63:0] GRF12_3_buffer [0:1];
  logic [63:0] GRF12_4_buffer [0:1];
  logic [63:0] GRF12_5_buffer [0:1];
  logic [63:0] GRF12_6_buffer [0:1];
  logic [63:0] GRF12_7_buffer [0:1];
  logic [63:0] GRF12_8_buffer [0:1];
  logic [63:0] GRF12_9_buffer [0:1];
  logic [63:0] GRF12_10_buffer [0:1];
  logic [63:0] GRF12_11_buffer [0:1];
  logic [63:0] GRF12_12_buffer [0:1];
  logic [63:0] GRF12_13_buffer [0:1];
  logic [63:0] GRF12_14_buffer [0:1];
  logic [63:0] GRF12_15_buffer [0:1];
  logic [63:0] GRF12_16_buffer [0:1];
  logic [63:0] GRF12_17_buffer [0:1];
  logic [63:0] GRF12_18_buffer [0:1];
  logic [63:0] GRF12_19_buffer [0:1];
  logic [63:0] GRF12_20_buffer [0:1];
  logic [63:0] GRF12_21_buffer [0:1];
  logic [63:0] GRF12_22_buffer [0:1];
  logic [63:0] GRF12_23_buffer [0:1];
  logic [63:0] GRF12_24_buffer [0:1];
  logic [63:0] GRF12_25_buffer [0:1];
  logic [63:0] GRF12_26_buffer [0:1];
  logic [63:0] GRF12_27_buffer [0:1];
  logic [63:0] GRF12_28_buffer [0:1];
  logic [63:0] GRF12_29_buffer [0:1];
  logic [63:0] GRF12_30_buffer [0:1];
  logic [63:0] GRF12_31_buffer [0:1];
  logic [63:0] GRF13_0_buffer [0:1];
  logic [63:0] GRF13_1_buffer [0:1];
  logic [63:0] GRF13_2_buffer [0:1];
  logic [63:0] GRF13_3_buffer [0:1];
  logic [63:0] GRF13_4_buffer [0:1];
  logic [63:0] GRF13_5_buffer [0:1];
  logic [63:0] GRF13_6_buffer [0:1];
  logic [63:0] GRF13_7_buffer [0:1];
  logic [63:0] GRF13_8_buffer [0:1];
  logic [63:0] GRF13_9_buffer [0:1];
  logic [63:0] GRF13_10_buffer [0:1];
  logic [63:0] GRF13_11_buffer [0:1];
  logic [63:0] GRF13_12_buffer [0:1];
  logic [63:0] GRF13_13_buffer [0:1];
  logic [63:0] GRF13_14_buffer [0:1];
  logic [63:0] GRF13_15_buffer [0:1];
  logic [63:0] GRF13_16_buffer [0:1];
  logic [63:0] GRF13_17_buffer [0:1];
  logic [63:0] GRF13_18_buffer [0:1];
  logic [63:0] GRF13_19_buffer [0:1];
  logic [63:0] GRF13_20_buffer [0:1];
  logic [63:0] GRF13_21_buffer [0:1];
  logic [63:0] GRF13_22_buffer [0:1];
  logic [63:0] GRF13_23_buffer [0:1];
  logic [63:0] GRF13_24_buffer [0:1];
  logic [63:0] GRF13_25_buffer [0:1];
  logic [63:0] GRF13_26_buffer [0:1];
  logic [63:0] GRF13_27_buffer [0:1];
  logic [63:0] GRF13_28_buffer [0:1];
  logic [63:0] GRF13_29_buffer [0:1];
  logic [63:0] GRF13_30_buffer [0:1];
  logic [63:0] GRF13_31_buffer [0:1];
  logic [63:0] GRF14_0_buffer [0:1];
  logic [63:0] GRF14_1_buffer [0:1];
  logic [63:0] GRF14_2_buffer [0:1];
  logic [63:0] GRF14_3_buffer [0:1];
  logic [63:0] GRF14_4_buffer [0:1];
  logic [63:0] GRF14_5_buffer [0:1];
  logic [63:0] GRF14_6_buffer [0:1];
  logic [63:0] GRF14_7_buffer [0:1];
  logic [63:0] GRF14_8_buffer [0:1];
  logic [63:0] GRF14_9_buffer [0:1];
  logic [63:0] GRF14_10_buffer [0:1];
  logic [63:0] GRF14_11_buffer [0:1];
  logic [63:0] GRF14_12_buffer [0:1];
  logic [63:0] GRF14_13_buffer [0:1];
  logic [63:0] GRF14_14_buffer [0:1];
  logic [63:0] GRF14_15_buffer [0:1];
  logic [63:0] GRF14_16_buffer [0:1];
  logic [63:0] GRF14_17_buffer [0:1];
  logic [63:0] GRF14_18_buffer [0:1];
  logic [63:0] GRF14_19_buffer [0:1];
  logic [63:0] GRF14_20_buffer [0:1];
  logic [63:0] GRF14_21_buffer [0:1];
  logic [63:0] GRF14_22_buffer [0:1];
  logic [63:0] GRF14_23_buffer [0:1];
  logic [63:0] GRF14_24_buffer [0:1];
  logic [63:0] GRF14_25_buffer [0:1];
  logic [63:0] GRF14_26_buffer [0:1];
  logic [63:0] GRF14_27_buffer [0:1];
  logic [63:0] GRF14_28_buffer [0:1];
  logic [63:0] GRF14_29_buffer [0:1];
  logic [63:0] GRF14_30_buffer [0:1];
  logic [63:0] GRF14_31_buffer [0:1];
  logic [63:0] GRF15_0_buffer [0:1];
  logic [63:0] GRF15_1_buffer [0:1];
  logic [63:0] GRF15_2_buffer [0:1];
  logic [63:0] GRF15_3_buffer [0:1];
  logic [63:0] GRF15_4_buffer [0:1];
  logic [63:0] GRF15_5_buffer [0:1];
  logic [63:0] GRF15_6_buffer [0:1];
  logic [63:0] GRF15_7_buffer [0:1];
  logic [63:0] GRF15_8_buffer [0:1];
  logic [63:0] GRF15_9_buffer [0:1];
  logic [63:0] GRF15_10_buffer [0:1];
  logic [63:0] GRF15_11_buffer [0:1];
  logic [63:0] GRF15_12_buffer [0:1];
  logic [63:0] GRF15_13_buffer [0:1];
  logic [63:0] GRF15_14_buffer [0:1];
  logic [63:0] GRF15_15_buffer [0:1];
  logic [63:0] GRF15_16_buffer [0:1];
  logic [63:0] GRF15_17_buffer [0:1];
  logic [63:0] GRF15_18_buffer [0:1];
  logic [63:0] GRF15_19_buffer [0:1];
  logic [63:0] GRF15_20_buffer [0:1];
  logic [63:0] GRF15_21_buffer [0:1];
  logic [63:0] GRF15_22_buffer [0:1];
  logic [63:0] GRF15_23_buffer [0:1];
  logic [63:0] GRF15_24_buffer [0:1];
  logic [63:0] GRF15_25_buffer [0:1];
  logic [63:0] GRF15_26_buffer [0:1];
  logic [63:0] GRF15_27_buffer [0:1];
  logic [63:0] GRF15_28_buffer [0:1];
  logic [63:0] GRF15_29_buffer [0:1];
  logic [63:0] GRF15_30_buffer [0:1];
  logic [63:0] GRF15_31_buffer [0:1];
  logic [63:0] GRF16_0_buffer [0:1];
  logic [63:0] GRF16_1_buffer [0:1];
  logic [63:0] GRF16_2_buffer [0:1];
  logic [63:0] GRF16_3_buffer [0:1];
  logic [63:0] GRF16_4_buffer [0:1];
  logic [63:0] GRF16_5_buffer [0:1];
  logic [63:0] GRF16_6_buffer [0:1];
  logic [63:0] GRF16_7_buffer [0:1];
  logic [63:0] GRF16_8_buffer [0:1];
  logic [63:0] GRF16_9_buffer [0:1];
  logic [63:0] GRF16_10_buffer [0:1];
  logic [63:0] GRF16_11_buffer [0:1];
  logic [63:0] GRF16_12_buffer [0:1];
  logic [63:0] GRF16_13_buffer [0:1];
  logic [63:0] GRF16_14_buffer [0:1];
  logic [63:0] GRF16_15_buffer [0:1];
  logic [63:0] GRF16_16_buffer [0:1];
  logic [63:0] GRF16_17_buffer [0:1];
  logic [63:0] GRF16_18_buffer [0:1];
  logic [63:0] GRF16_19_buffer [0:1];
  logic [63:0] GRF16_20_buffer [0:1];
  logic [63:0] GRF16_21_buffer [0:1];
  logic [63:0] GRF16_22_buffer [0:1];
  logic [63:0] GRF16_23_buffer [0:1];
  logic [63:0] GRF16_24_buffer [0:1];
  logic [63:0] GRF16_25_buffer [0:1];
  logic [63:0] GRF16_26_buffer [0:1];
  logic [63:0] GRF16_27_buffer [0:1];
  logic [63:0] GRF16_28_buffer [0:1];
  logic [63:0] GRF16_29_buffer [0:1];
  logic [63:0] GRF16_30_buffer [0:1];
  logic [63:0] GRF16_31_buffer [0:1];
  logic [63:0] GRF17_0_buffer [0:1];
  logic [63:0] GRF17_1_buffer [0:1];
  logic [63:0] GRF17_2_buffer [0:1];
  logic [63:0] GRF17_3_buffer [0:1];
  logic [63:0] GRF17_4_buffer [0:1];
  logic [63:0] GRF17_5_buffer [0:1];
  logic [63:0] GRF17_6_buffer [0:1];
  logic [63:0] GRF17_7_buffer [0:1];
  logic [63:0] GRF17_8_buffer [0:1];
  logic [63:0] GRF17_9_buffer [0:1];
  logic [63:0] GRF17_10_buffer [0:1];
  logic [63:0] GRF17_11_buffer [0:1];
  logic [63:0] GRF17_12_buffer [0:1];
  logic [63:0] GRF17_13_buffer [0:1];
  logic [63:0] GRF17_14_buffer [0:1];
  logic [63:0] GRF17_15_buffer [0:1];
  logic [63:0] GRF17_16_buffer [0:1];
  logic [63:0] GRF17_17_buffer [0:1];
  logic [63:0] GRF17_18_buffer [0:1];
  logic [63:0] GRF17_19_buffer [0:1];
  logic [63:0] GRF17_20_buffer [0:1];
  logic [63:0] GRF17_21_buffer [0:1];
  logic [63:0] GRF17_22_buffer [0:1];
  logic [63:0] GRF17_23_buffer [0:1];
  logic [63:0] GRF17_24_buffer [0:1];
  logic [63:0] GRF17_25_buffer [0:1];
  logic [63:0] GRF17_26_buffer [0:1];
  logic [63:0] GRF17_27_buffer [0:1];
  logic [63:0] GRF17_28_buffer [0:1];
  logic [63:0] GRF17_29_buffer [0:1];
  logic [63:0] GRF17_30_buffer [0:1];
  logic [63:0] GRF17_31_buffer [0:1];
  logic [63:0] GRF18_0_buffer [0:1];
  logic [63:0] GRF18_1_buffer [0:1];
  logic [63:0] GRF18_2_buffer [0:1];
  logic [63:0] GRF18_3_buffer [0:1];
  logic [63:0] GRF18_4_buffer [0:1];
  logic [63:0] GRF18_5_buffer [0:1];
  logic [63:0] GRF18_6_buffer [0:1];
  logic [63:0] GRF18_7_buffer [0:1];
  logic [63:0] GRF18_8_buffer [0:1];
  logic [63:0] GRF18_9_buffer [0:1];
  logic [63:0] GRF18_10_buffer [0:1];
  logic [63:0] GRF18_11_buffer [0:1];
  logic [63:0] GRF18_12_buffer [0:1];
  logic [63:0] GRF18_13_buffer [0:1];
  logic [63:0] GRF18_14_buffer [0:1];
  logic [63:0] GRF18_15_buffer [0:1];
  logic [63:0] GRF18_16_buffer [0:1];
  logic [63:0] GRF18_17_buffer [0:1];
  logic [63:0] GRF18_18_buffer [0:1];
  logic [63:0] GRF18_19_buffer [0:1];
  logic [63:0] GRF18_20_buffer [0:1];
  logic [63:0] GRF18_21_buffer [0:1];
  logic [63:0] GRF18_22_buffer [0:1];
  logic [63:0] GRF18_23_buffer [0:1];
  logic [63:0] GRF18_24_buffer [0:1];
  logic [63:0] GRF18_25_buffer [0:1];
  logic [63:0] GRF18_26_buffer [0:1];
  logic [63:0] GRF18_27_buffer [0:1];
  logic [63:0] GRF18_28_buffer [0:1];
  logic [63:0] GRF18_29_buffer [0:1];
  logic [63:0] GRF18_30_buffer [0:1];
  logic [63:0] GRF18_31_buffer [0:1];
  logic [63:0] GRF19_0_buffer [0:1];
  logic [63:0] GRF19_1_buffer [0:1];
  logic [63:0] GRF19_2_buffer [0:1];
  logic [63:0] GRF19_3_buffer [0:1];
  logic [63:0] GRF19_4_buffer [0:1];
  logic [63:0] GRF19_5_buffer [0:1];
  logic [63:0] GRF19_6_buffer [0:1];
  logic [63:0] GRF19_7_buffer [0:1];
  logic [63:0] GRF19_8_buffer [0:1];
  logic [63:0] GRF19_9_buffer [0:1];
  logic [63:0] GRF19_10_buffer [0:1];
  logic [63:0] GRF19_11_buffer [0:1];
  logic [63:0] GRF19_12_buffer [0:1];
  logic [63:0] GRF19_13_buffer [0:1];
  logic [63:0] GRF19_14_buffer [0:1];
  logic [63:0] GRF19_15_buffer [0:1];
  logic [63:0] GRF19_16_buffer [0:1];
  logic [63:0] GRF19_17_buffer [0:1];
  logic [63:0] GRF19_18_buffer [0:1];
  logic [63:0] GRF19_19_buffer [0:1];
  logic [63:0] GRF19_20_buffer [0:1];
  logic [63:0] GRF19_21_buffer [0:1];
  logic [63:0] GRF19_22_buffer [0:1];
  logic [63:0] GRF19_23_buffer [0:1];
  logic [63:0] GRF19_24_buffer [0:1];
  logic [63:0] GRF19_25_buffer [0:1];
  logic [63:0] GRF19_26_buffer [0:1];
  logic [63:0] GRF19_27_buffer [0:1];
  logic [63:0] GRF19_28_buffer [0:1];
  logic [63:0] GRF19_29_buffer [0:1];
  logic [63:0] GRF19_30_buffer [0:1];
  logic [63:0] GRF19_31_buffer [0:1];
  logic [63:0] GRF20_0_buffer [0:1];
  logic [63:0] GRF20_1_buffer [0:1];
  logic [63:0] GRF20_2_buffer [0:1];
  logic [63:0] GRF20_3_buffer [0:1];
  logic [63:0] GRF20_4_buffer [0:1];
  logic [63:0] GRF20_5_buffer [0:1];
  logic [63:0] GRF20_6_buffer [0:1];
  logic [63:0] GRF20_7_buffer [0:1];
  logic [63:0] GRF20_8_buffer [0:1];
  logic [63:0] GRF20_9_buffer [0:1];
  logic [63:0] GRF20_10_buffer [0:1];
  logic [63:0] GRF20_11_buffer [0:1];
  logic [63:0] GRF20_12_buffer [0:1];
  logic [63:0] GRF20_13_buffer [0:1];
  logic [63:0] GRF20_14_buffer [0:1];
  logic [63:0] GRF20_15_buffer [0:1];
  logic [63:0] GRF20_16_buffer [0:1];
  logic [63:0] GRF20_17_buffer [0:1];
  logic [63:0] GRF20_18_buffer [0:1];
  logic [63:0] GRF20_19_buffer [0:1];
  logic [63:0] GRF20_20_buffer [0:1];
  logic [63:0] GRF20_21_buffer [0:1];
  logic [63:0] GRF20_22_buffer [0:1];
  logic [63:0] GRF20_23_buffer [0:1];
  logic [63:0] GRF20_24_buffer [0:1];
  logic [63:0] GRF20_25_buffer [0:1];
  logic [63:0] GRF20_26_buffer [0:1];
  logic [63:0] GRF20_27_buffer [0:1];
  logic [63:0] GRF20_28_buffer [0:1];
  logic [63:0] GRF20_29_buffer [0:1];
  logic [63:0] GRF20_30_buffer [0:1];
  logic [63:0] GRF20_31_buffer [0:1];
  logic [63:0] GRF21_0_buffer [0:1];
  logic [63:0] GRF21_1_buffer [0:1];
  logic [63:0] GRF21_2_buffer [0:1];
  logic [63:0] GRF21_3_buffer [0:1];
  logic [63:0] GRF21_4_buffer [0:1];
  logic [63:0] GRF21_5_buffer [0:1];
  logic [63:0] GRF21_6_buffer [0:1];
  logic [63:0] GRF21_7_buffer [0:1];
  logic [63:0] GRF21_8_buffer [0:1];
  logic [63:0] GRF21_9_buffer [0:1];
  logic [63:0] GRF21_10_buffer [0:1];
  logic [63:0] GRF21_11_buffer [0:1];
  logic [63:0] GRF21_12_buffer [0:1];
  logic [63:0] GRF21_13_buffer [0:1];
  logic [63:0] GRF21_14_buffer [0:1];
  logic [63:0] GRF21_15_buffer [0:1];
  logic [63:0] GRF21_16_buffer [0:1];
  logic [63:0] GRF21_17_buffer [0:1];
  logic [63:0] GRF21_18_buffer [0:1];
  logic [63:0] GRF21_19_buffer [0:1];
  logic [63:0] GRF21_20_buffer [0:1];
  logic [63:0] GRF21_21_buffer [0:1];
  logic [63:0] GRF21_22_buffer [0:1];
  logic [63:0] GRF21_23_buffer [0:1];
  logic [63:0] GRF21_24_buffer [0:1];
  logic [63:0] GRF21_25_buffer [0:1];
  logic [63:0] GRF21_26_buffer [0:1];
  logic [63:0] GRF21_27_buffer [0:1];
  logic [63:0] GRF21_28_buffer [0:1];
  logic [63:0] GRF21_29_buffer [0:1];
  logic [63:0] GRF21_30_buffer [0:1];
  logic [63:0] GRF21_31_buffer [0:1];
  logic [63:0] GRF22_0_buffer [0:1];
  logic [63:0] GRF22_1_buffer [0:1];
  logic [63:0] GRF22_2_buffer [0:1];
  logic [63:0] GRF22_3_buffer [0:1];
  logic [63:0] GRF22_4_buffer [0:1];
  logic [63:0] GRF22_5_buffer [0:1];
  logic [63:0] GRF22_6_buffer [0:1];
  logic [63:0] GRF22_7_buffer [0:1];
  logic [63:0] GRF22_8_buffer [0:1];
  logic [63:0] GRF22_9_buffer [0:1];
  logic [63:0] GRF22_10_buffer [0:1];
  logic [63:0] GRF22_11_buffer [0:1];
  logic [63:0] GRF22_12_buffer [0:1];
  logic [63:0] GRF22_13_buffer [0:1];
  logic [63:0] GRF22_14_buffer [0:1];
  logic [63:0] GRF22_15_buffer [0:1];
  logic [63:0] GRF22_16_buffer [0:1];
  logic [63:0] GRF22_17_buffer [0:1];
  logic [63:0] GRF22_18_buffer [0:1];
  logic [63:0] GRF22_19_buffer [0:1];
  logic [63:0] GRF22_20_buffer [0:1];
  logic [63:0] GRF22_21_buffer [0:1];
  logic [63:0] GRF22_22_buffer [0:1];
  logic [63:0] GRF22_23_buffer [0:1];
  logic [63:0] GRF22_24_buffer [0:1];
  logic [63:0] GRF22_25_buffer [0:1];
  logic [63:0] GRF22_26_buffer [0:1];
  logic [63:0] GRF22_27_buffer [0:1];
  logic [63:0] GRF22_28_buffer [0:1];
  logic [63:0] GRF22_29_buffer [0:1];
  logic [63:0] GRF22_30_buffer [0:1];
  logic [63:0] GRF22_31_buffer [0:1];
  logic [63:0] GRF23_0_buffer [0:1];
  logic [63:0] GRF23_1_buffer [0:1];
  logic [63:0] GRF23_2_buffer [0:1];
  logic [63:0] GRF23_3_buffer [0:1];
  logic [63:0] GRF23_4_buffer [0:1];
  logic [63:0] GRF23_5_buffer [0:1];
  logic [63:0] GRF23_6_buffer [0:1];
  logic [63:0] GRF23_7_buffer [0:1];
  logic [63:0] GRF23_8_buffer [0:1];
  logic [63:0] GRF23_9_buffer [0:1];
  logic [63:0] GRF23_10_buffer [0:1];
  logic [63:0] GRF23_11_buffer [0:1];
  logic [63:0] GRF23_12_buffer [0:1];
  logic [63:0] GRF23_13_buffer [0:1];
  logic [63:0] GRF23_14_buffer [0:1];
  logic [63:0] GRF23_15_buffer [0:1];
  logic [63:0] GRF23_16_buffer [0:1];
  logic [63:0] GRF23_17_buffer [0:1];
  logic [63:0] GRF23_18_buffer [0:1];
  logic [63:0] GRF23_19_buffer [0:1];
  logic [63:0] GRF23_20_buffer [0:1];
  logic [63:0] GRF23_21_buffer [0:1];
  logic [63:0] GRF23_22_buffer [0:1];
  logic [63:0] GRF23_23_buffer [0:1];
  logic [63:0] GRF23_24_buffer [0:1];
  logic [63:0] GRF23_25_buffer [0:1];
  logic [63:0] GRF23_26_buffer [0:1];
  logic [63:0] GRF23_27_buffer [0:1];
  logic [63:0] GRF23_28_buffer [0:1];
  logic [63:0] GRF23_29_buffer [0:1];
  logic [63:0] GRF23_30_buffer [0:1];
  logic [63:0] GRF23_31_buffer [0:1];
  logic [63:0] GRF24_0_buffer [0:1];
  logic [63:0] GRF24_1_buffer [0:1];
  logic [63:0] GRF24_2_buffer [0:1];
  logic [63:0] GRF24_3_buffer [0:1];
  logic [63:0] GRF24_4_buffer [0:1];
  logic [63:0] GRF24_5_buffer [0:1];
  logic [63:0] GRF24_6_buffer [0:1];
  logic [63:0] GRF24_7_buffer [0:1];
  logic [63:0] GRF24_8_buffer [0:1];
  logic [63:0] GRF24_9_buffer [0:1];
  logic [63:0] GRF24_10_buffer [0:1];
  logic [63:0] GRF24_11_buffer [0:1];
  logic [63:0] GRF24_12_buffer [0:1];
  logic [63:0] GRF24_13_buffer [0:1];
  logic [63:0] GRF24_14_buffer [0:1];
  logic [63:0] GRF24_15_buffer [0:1];
  logic [63:0] GRF24_16_buffer [0:1];
  logic [63:0] GRF24_17_buffer [0:1];
  logic [63:0] GRF24_18_buffer [0:1];
  logic [63:0] GRF24_19_buffer [0:1];
  logic [63:0] GRF24_20_buffer [0:1];
  logic [63:0] GRF24_21_buffer [0:1];
  logic [63:0] GRF24_22_buffer [0:1];
  logic [63:0] GRF24_23_buffer [0:1];
  logic [63:0] GRF24_24_buffer [0:1];
  logic [63:0] GRF24_25_buffer [0:1];
  logic [63:0] GRF24_26_buffer [0:1];
  logic [63:0] GRF24_27_buffer [0:1];
  logic [63:0] GRF24_28_buffer [0:1];
  logic [63:0] GRF24_29_buffer [0:1];
  logic [63:0] GRF24_30_buffer [0:1];
  logic [63:0] GRF24_31_buffer [0:1];
  logic [63:0] GRF25_0_buffer [0:1];
  logic [63:0] GRF25_1_buffer [0:1];
  logic [63:0] GRF25_2_buffer [0:1];
  logic [63:0] GRF25_3_buffer [0:1];
  logic [63:0] GRF25_4_buffer [0:1];
  logic [63:0] GRF25_5_buffer [0:1];
  logic [63:0] GRF25_6_buffer [0:1];
  logic [63:0] GRF25_7_buffer [0:1];
  logic [63:0] GRF25_8_buffer [0:1];
  logic [63:0] GRF25_9_buffer [0:1];
  logic [63:0] GRF25_10_buffer [0:1];
  logic [63:0] GRF25_11_buffer [0:1];
  logic [63:0] GRF25_12_buffer [0:1];
  logic [63:0] GRF25_13_buffer [0:1];
  logic [63:0] GRF25_14_buffer [0:1];
  logic [63:0] GRF25_15_buffer [0:1];
  logic [63:0] GRF25_16_buffer [0:1];
  logic [63:0] GRF25_17_buffer [0:1];
  logic [63:0] GRF25_18_buffer [0:1];
  logic [63:0] GRF25_19_buffer [0:1];
  logic [63:0] GRF25_20_buffer [0:1];
  logic [63:0] GRF25_21_buffer [0:1];
  logic [63:0] GRF25_22_buffer [0:1];
  logic [63:0] GRF25_23_buffer [0:1];
  logic [63:0] GRF25_24_buffer [0:1];
  logic [63:0] GRF25_25_buffer [0:1];
  logic [63:0] GRF25_26_buffer [0:1];
  logic [63:0] GRF25_27_buffer [0:1];
  logic [63:0] GRF25_28_buffer [0:1];
  logic [63:0] GRF25_29_buffer [0:1];
  logic [63:0] GRF25_30_buffer [0:1];
  logic [63:0] GRF25_31_buffer [0:1];
  logic [63:0] GRF26_0_buffer [0:1];
  logic [63:0] GRF26_1_buffer [0:1];
  logic [63:0] GRF26_2_buffer [0:1];
  logic [63:0] GRF26_3_buffer [0:1];
  logic [63:0] GRF26_4_buffer [0:1];
  logic [63:0] GRF26_5_buffer [0:1];
  logic [63:0] GRF26_6_buffer [0:1];
  logic [63:0] GRF26_7_buffer [0:1];
  logic [63:0] GRF26_8_buffer [0:1];
  logic [63:0] GRF26_9_buffer [0:1];
  logic [63:0] GRF26_10_buffer [0:1];
  logic [63:0] GRF26_11_buffer [0:1];
  logic [63:0] GRF26_12_buffer [0:1];
  logic [63:0] GRF26_13_buffer [0:1];
  logic [63:0] GRF26_14_buffer [0:1];
  logic [63:0] GRF26_15_buffer [0:1];
  logic [63:0] GRF26_16_buffer [0:1];
  logic [63:0] GRF26_17_buffer [0:1];
  logic [63:0] GRF26_18_buffer [0:1];
  logic [63:0] GRF26_19_buffer [0:1];
  logic [63:0] GRF26_20_buffer [0:1];
  logic [63:0] GRF26_21_buffer [0:1];
  logic [63:0] GRF26_22_buffer [0:1];
  logic [63:0] GRF26_23_buffer [0:1];
  logic [63:0] GRF26_24_buffer [0:1];
  logic [63:0] GRF26_25_buffer [0:1];
  logic [63:0] GRF26_26_buffer [0:1];
  logic [63:0] GRF26_27_buffer [0:1];
  logic [63:0] GRF26_28_buffer [0:1];
  logic [63:0] GRF26_29_buffer [0:1];
  logic [63:0] GRF26_30_buffer [0:1];
  logic [63:0] GRF26_31_buffer [0:1];
  logic [63:0] GRF27_0_buffer [0:1];
  logic [63:0] GRF27_1_buffer [0:1];
  logic [63:0] GRF27_2_buffer [0:1];
  logic [63:0] GRF27_3_buffer [0:1];
  logic [63:0] GRF27_4_buffer [0:1];
  logic [63:0] GRF27_5_buffer [0:1];
  logic [63:0] GRF27_6_buffer [0:1];
  logic [63:0] GRF27_7_buffer [0:1];
  logic [63:0] GRF27_8_buffer [0:1];
  logic [63:0] GRF27_9_buffer [0:1];
  logic [63:0] GRF27_10_buffer [0:1];
  logic [63:0] GRF27_11_buffer [0:1];
  logic [63:0] GRF27_12_buffer [0:1];
  logic [63:0] GRF27_13_buffer [0:1];
  logic [63:0] GRF27_14_buffer [0:1];
  logic [63:0] GRF27_15_buffer [0:1];
  logic [63:0] GRF27_16_buffer [0:1];
  logic [63:0] GRF27_17_buffer [0:1];
  logic [63:0] GRF27_18_buffer [0:1];
  logic [63:0] GRF27_19_buffer [0:1];
  logic [63:0] GRF27_20_buffer [0:1];
  logic [63:0] GRF27_21_buffer [0:1];
  logic [63:0] GRF27_22_buffer [0:1];
  logic [63:0] GRF27_23_buffer [0:1];
  logic [63:0] GRF27_24_buffer [0:1];
  logic [63:0] GRF27_25_buffer [0:1];
  logic [63:0] GRF27_26_buffer [0:1];
  logic [63:0] GRF27_27_buffer [0:1];
  logic [63:0] GRF27_28_buffer [0:1];
  logic [63:0] GRF27_29_buffer [0:1];
  logic [63:0] GRF27_30_buffer [0:1];
  logic [63:0] GRF27_31_buffer [0:1];
  logic [63:0] GRF28_0_buffer [0:1];
  logic [63:0] GRF28_1_buffer [0:1];
  logic [63:0] GRF28_2_buffer [0:1];
  logic [63:0] GRF28_3_buffer [0:1];
  logic [63:0] GRF28_4_buffer [0:1];
  logic [63:0] GRF28_5_buffer [0:1];
  logic [63:0] GRF28_6_buffer [0:1];
  logic [63:0] GRF28_7_buffer [0:1];
  logic [63:0] GRF28_8_buffer [0:1];
  logic [63:0] GRF28_9_buffer [0:1];
  logic [63:0] GRF28_10_buffer [0:1];
  logic [63:0] GRF28_11_buffer [0:1];
  logic [63:0] GRF28_12_buffer [0:1];
  logic [63:0] GRF28_13_buffer [0:1];
  logic [63:0] GRF28_14_buffer [0:1];
  logic [63:0] GRF28_15_buffer [0:1];
  logic [63:0] GRF28_16_buffer [0:1];
  logic [63:0] GRF28_17_buffer [0:1];
  logic [63:0] GRF28_18_buffer [0:1];
  logic [63:0] GRF28_19_buffer [0:1];
  logic [63:0] GRF28_20_buffer [0:1];
  logic [63:0] GRF28_21_buffer [0:1];
  logic [63:0] GRF28_22_buffer [0:1];
  logic [63:0] GRF28_23_buffer [0:1];
  logic [63:0] GRF28_24_buffer [0:1];
  logic [63:0] GRF28_25_buffer [0:1];
  logic [63:0] GRF28_26_buffer [0:1];
  logic [63:0] GRF28_27_buffer [0:1];
  logic [63:0] GRF28_28_buffer [0:1];
  logic [63:0] GRF28_29_buffer [0:1];
  logic [63:0] GRF28_30_buffer [0:1];
  logic [63:0] GRF28_31_buffer [0:1];
  logic [63:0] GRF29_0_buffer [0:1];
  logic [63:0] GRF29_1_buffer [0:1];
  logic [63:0] GRF29_2_buffer [0:1];
  logic [63:0] GRF29_3_buffer [0:1];
  logic [63:0] GRF29_4_buffer [0:1];
  logic [63:0] GRF29_5_buffer [0:1];
  logic [63:0] GRF29_6_buffer [0:1];
  logic [63:0] GRF29_7_buffer [0:1];
  logic [63:0] GRF29_8_buffer [0:1];
  logic [63:0] GRF29_9_buffer [0:1];
  logic [63:0] GRF29_10_buffer [0:1];
  logic [63:0] GRF29_11_buffer [0:1];
  logic [63:0] GRF29_12_buffer [0:1];
  logic [63:0] GRF29_13_buffer [0:1];
  logic [63:0] GRF29_14_buffer [0:1];
  logic [63:0] GRF29_15_buffer [0:1];
  logic [63:0] GRF29_16_buffer [0:1];
  logic [63:0] GRF29_17_buffer [0:1];
  logic [63:0] GRF29_18_buffer [0:1];
  logic [63:0] GRF29_19_buffer [0:1];
  logic [63:0] GRF29_20_buffer [0:1];
  logic [63:0] GRF29_21_buffer [0:1];
  logic [63:0] GRF29_22_buffer [0:1];
  logic [63:0] GRF29_23_buffer [0:1];
  logic [63:0] GRF29_24_buffer [0:1];
  logic [63:0] GRF29_25_buffer [0:1];
  logic [63:0] GRF29_26_buffer [0:1];
  logic [63:0] GRF29_27_buffer [0:1];
  logic [63:0] GRF29_28_buffer [0:1];
  logic [63:0] GRF29_29_buffer [0:1];
  logic [63:0] GRF29_30_buffer [0:1];
  logic [63:0] GRF29_31_buffer [0:1];
  logic [63:0] GRF30_0_buffer [0:1];
  logic [63:0] GRF30_1_buffer [0:1];
  logic [63:0] GRF30_2_buffer [0:1];
  logic [63:0] GRF30_3_buffer [0:1];
  logic [63:0] GRF30_4_buffer [0:1];
  logic [63:0] GRF30_5_buffer [0:1];
  logic [63:0] GRF30_6_buffer [0:1];
  logic [63:0] GRF30_7_buffer [0:1];
  logic [63:0] GRF30_8_buffer [0:1];
  logic [63:0] GRF30_9_buffer [0:1];
  logic [63:0] GRF30_10_buffer [0:1];
  logic [63:0] GRF30_11_buffer [0:1];
  logic [63:0] GRF30_12_buffer [0:1];
  logic [63:0] GRF30_13_buffer [0:1];
  logic [63:0] GRF30_14_buffer [0:1];
  logic [63:0] GRF30_15_buffer [0:1];
  logic [63:0] GRF30_16_buffer [0:1];
  logic [63:0] GRF30_17_buffer [0:1];
  logic [63:0] GRF30_18_buffer [0:1];
  logic [63:0] GRF30_19_buffer [0:1];
  logic [63:0] GRF30_20_buffer [0:1];
  logic [63:0] GRF30_21_buffer [0:1];
  logic [63:0] GRF30_22_buffer [0:1];
  logic [63:0] GRF30_23_buffer [0:1];
  logic [63:0] GRF30_24_buffer [0:1];
  logic [63:0] GRF30_25_buffer [0:1];
  logic [63:0] GRF30_26_buffer [0:1];
  logic [63:0] GRF30_27_buffer [0:1];
  logic [63:0] GRF30_28_buffer [0:1];
  logic [63:0] GRF30_29_buffer [0:1];
  logic [63:0] GRF30_30_buffer [0:1];
  logic [63:0] GRF30_31_buffer [0:1];
  logic [63:0] GRF31_0_buffer [0:1];
  logic [63:0] GRF31_1_buffer [0:1];
  logic [63:0] GRF31_2_buffer [0:1];
  logic [63:0] GRF31_3_buffer [0:1];
  logic [63:0] GRF31_4_buffer [0:1];
  logic [63:0] GRF31_5_buffer [0:1];
  logic [63:0] GRF31_6_buffer [0:1];
  logic [63:0] GRF31_7_buffer [0:1];
  logic [63:0] GRF31_8_buffer [0:1];
  logic [63:0] GRF31_9_buffer [0:1];
  logic [63:0] GRF31_10_buffer [0:1];
  logic [63:0] GRF31_11_buffer [0:1];
  logic [63:0] GRF31_12_buffer [0:1];
  logic [63:0] GRF31_13_buffer [0:1];
  logic [63:0] GRF31_14_buffer [0:1];
  logic [63:0] GRF31_15_buffer [0:1];
  logic [63:0] GRF31_16_buffer [0:1];
  logic [63:0] GRF31_17_buffer [0:1];
  logic [63:0] GRF31_18_buffer [0:1];
  logic [63:0] GRF31_19_buffer [0:1];
  logic [63:0] GRF31_20_buffer [0:1];
  logic [63:0] GRF31_21_buffer [0:1];
  logic [63:0] GRF31_22_buffer [0:1];
  logic [63:0] GRF31_23_buffer [0:1];
  logic [63:0] GRF31_24_buffer [0:1];
  logic [63:0] GRF31_25_buffer [0:1];
  logic [63:0] GRF31_26_buffer [0:1];
  logic [63:0] GRF31_27_buffer [0:1];
  logic [63:0] GRF31_28_buffer [0:1];
  logic [63:0] GRF31_29_buffer [0:1];
  logic [63:0] GRF31_30_buffer [0:1];
  logic [63:0] GRF31_31_buffer [0:1];
  logic [63:0] GRF32_0_buffer [0:1];
  logic [63:0] GRF32_1_buffer [0:1];
  logic [63:0] GRF32_2_buffer [0:1];
  logic [63:0] GRF32_3_buffer [0:1];
  logic [63:0] GRF32_4_buffer [0:1];
  logic [63:0] GRF32_5_buffer [0:1];
  logic [63:0] GRF32_6_buffer [0:1];
  logic [63:0] GRF32_7_buffer [0:1];
  logic [63:0] GRF32_8_buffer [0:1];
  logic [63:0] GRF32_9_buffer [0:1];
  logic [63:0] GRF32_10_buffer [0:1];
  logic [63:0] GRF32_11_buffer [0:1];
  logic [63:0] GRF32_12_buffer [0:1];
  logic [63:0] GRF32_13_buffer [0:1];
  logic [63:0] GRF32_14_buffer [0:1];
  logic [63:0] GRF32_15_buffer [0:1];
  logic [63:0] GRF32_16_buffer [0:1];
  logic [63:0] GRF32_17_buffer [0:1];
  logic [63:0] GRF32_18_buffer [0:1];
  logic [63:0] GRF32_19_buffer [0:1];
  logic [63:0] GRF32_20_buffer [0:1];
  logic [63:0] GRF32_21_buffer [0:1];
  logic [63:0] GRF32_22_buffer [0:1];
  logic [63:0] GRF32_23_buffer [0:1];
  logic [63:0] GRF32_24_buffer [0:1];
  logic [63:0] GRF32_25_buffer [0:1];
  logic [63:0] GRF32_26_buffer [0:1];
  logic [63:0] GRF32_27_buffer [0:1];
  logic [63:0] GRF32_28_buffer [0:1];
  logic [63:0] GRF32_29_buffer [0:1];
  logic [63:0] GRF32_30_buffer [0:1];
  logic [63:0] GRF32_31_buffer [0:1];
  logic [63:0] GRF33_0_buffer [0:1];
  logic [63:0] GRF33_1_buffer [0:1];
  logic [63:0] GRF33_2_buffer [0:1];
  logic [63:0] GRF33_3_buffer [0:1];
  logic [63:0] GRF33_4_buffer [0:1];
  logic [63:0] GRF33_5_buffer [0:1];
  logic [63:0] GRF33_6_buffer [0:1];
  logic [63:0] GRF33_7_buffer [0:1];
  logic [63:0] GRF33_8_buffer [0:1];
  logic [63:0] GRF33_9_buffer [0:1];
  logic [63:0] GRF33_10_buffer [0:1];
  logic [63:0] GRF33_11_buffer [0:1];
  logic [63:0] GRF33_12_buffer [0:1];
  logic [63:0] GRF33_13_buffer [0:1];
  logic [63:0] GRF33_14_buffer [0:1];
  logic [63:0] GRF33_15_buffer [0:1];
  logic [63:0] GRF33_16_buffer [0:1];
  logic [63:0] GRF33_17_buffer [0:1];
  logic [63:0] GRF33_18_buffer [0:1];
  logic [63:0] GRF33_19_buffer [0:1];
  logic [63:0] GRF33_20_buffer [0:1];
  logic [63:0] GRF33_21_buffer [0:1];
  logic [63:0] GRF33_22_buffer [0:1];
  logic [63:0] GRF33_23_buffer [0:1];
  logic [63:0] GRF33_24_buffer [0:1];
  logic [63:0] GRF33_25_buffer [0:1];
  logic [63:0] GRF33_26_buffer [0:1];
  logic [63:0] GRF33_27_buffer [0:1];
  logic [63:0] GRF33_28_buffer [0:1];
  logic [63:0] GRF33_29_buffer [0:1];
  logic [63:0] GRF33_30_buffer [0:1];
  logic [63:0] GRF33_31_buffer [0:1];
  logic [63:0] GRF34_0_buffer [0:1];
  logic [63:0] GRF34_1_buffer [0:1];
  logic [63:0] GRF34_2_buffer [0:1];
  logic [63:0] GRF34_3_buffer [0:1];
  logic [63:0] GRF34_4_buffer [0:1];
  logic [63:0] GRF34_5_buffer [0:1];
  logic [63:0] GRF34_6_buffer [0:1];
  logic [63:0] GRF34_7_buffer [0:1];
  logic [63:0] GRF34_8_buffer [0:1];
  logic [63:0] GRF34_9_buffer [0:1];
  logic [63:0] GRF34_10_buffer [0:1];
  logic [63:0] GRF34_11_buffer [0:1];
  logic [63:0] GRF34_12_buffer [0:1];
  logic [63:0] GRF34_13_buffer [0:1];
  logic [63:0] GRF34_14_buffer [0:1];
  logic [63:0] GRF34_15_buffer [0:1];
  logic [63:0] GRF34_16_buffer [0:1];
  logic [63:0] GRF34_17_buffer [0:1];
  logic [63:0] GRF34_18_buffer [0:1];
  logic [63:0] GRF34_19_buffer [0:1];
  logic [63:0] GRF34_20_buffer [0:1];
  logic [63:0] GRF34_21_buffer [0:1];
  logic [63:0] GRF34_22_buffer [0:1];
  logic [63:0] GRF34_23_buffer [0:1];
  logic [63:0] GRF34_24_buffer [0:1];
  logic [63:0] GRF34_25_buffer [0:1];
  logic [63:0] GRF34_26_buffer [0:1];
  logic [63:0] GRF34_27_buffer [0:1];
  logic [63:0] GRF34_28_buffer [0:1];
  logic [63:0] GRF34_29_buffer [0:1];
  logic [63:0] GRF34_30_buffer [0:1];
  logic [63:0] GRF34_31_buffer [0:1];
  logic [63:0] GRF35_0_buffer [0:1];
  logic [63:0] GRF35_1_buffer [0:1];
  logic [63:0] GRF35_2_buffer [0:1];
  logic [63:0] GRF35_3_buffer [0:1];
  logic [63:0] GRF35_4_buffer [0:1];
  logic [63:0] GRF35_5_buffer [0:1];
  logic [63:0] GRF35_6_buffer [0:1];
  logic [63:0] GRF35_7_buffer [0:1];
  logic [63:0] GRF35_8_buffer [0:1];
  logic [63:0] GRF35_9_buffer [0:1];
  logic [63:0] GRF35_10_buffer [0:1];
  logic [63:0] GRF35_11_buffer [0:1];
  logic [63:0] GRF35_12_buffer [0:1];
  logic [63:0] GRF35_13_buffer [0:1];
  logic [63:0] GRF35_14_buffer [0:1];
  logic [63:0] GRF35_15_buffer [0:1];
  logic [63:0] GRF35_16_buffer [0:1];
  logic [63:0] GRF35_17_buffer [0:1];
  logic [63:0] GRF35_18_buffer [0:1];
  logic [63:0] GRF35_19_buffer [0:1];
  logic [63:0] GRF35_20_buffer [0:1];
  logic [63:0] GRF35_21_buffer [0:1];
  logic [63:0] GRF35_22_buffer [0:1];
  logic [63:0] GRF35_23_buffer [0:1];
  logic [63:0] GRF35_24_buffer [0:1];
  logic [63:0] GRF35_25_buffer [0:1];
  logic [63:0] GRF35_26_buffer [0:1];
  logic [63:0] GRF35_27_buffer [0:1];
  logic [63:0] GRF35_28_buffer [0:1];
  logic [63:0] GRF35_29_buffer [0:1];
  logic [63:0] GRF35_30_buffer [0:1];
  logic [63:0] GRF35_31_buffer [0:1];
  logic [63:0] GRF36_0_buffer [0:1];
  logic [63:0] GRF36_1_buffer [0:1];
  logic [63:0] GRF36_2_buffer [0:1];
  logic [63:0] GRF36_3_buffer [0:1];
  logic [63:0] GRF36_4_buffer [0:1];
  logic [63:0] GRF36_5_buffer [0:1];
  logic [63:0] GRF36_6_buffer [0:1];
  logic [63:0] GRF36_7_buffer [0:1];
  logic [63:0] GRF36_8_buffer [0:1];
  logic [63:0] GRF36_9_buffer [0:1];
  logic [63:0] GRF36_10_buffer [0:1];
  logic [63:0] GRF36_11_buffer [0:1];
  logic [63:0] GRF36_12_buffer [0:1];
  logic [63:0] GRF36_13_buffer [0:1];
  logic [63:0] GRF36_14_buffer [0:1];
  logic [63:0] GRF36_15_buffer [0:1];
  logic [63:0] GRF36_16_buffer [0:1];
  logic [63:0] GRF36_17_buffer [0:1];
  logic [63:0] GRF36_18_buffer [0:1];
  logic [63:0] GRF36_19_buffer [0:1];
  logic [63:0] GRF36_20_buffer [0:1];
  logic [63:0] GRF36_21_buffer [0:1];
  logic [63:0] GRF36_22_buffer [0:1];
  logic [63:0] GRF36_23_buffer [0:1];
  logic [63:0] GRF36_24_buffer [0:1];
  logic [63:0] GRF36_25_buffer [0:1];
  logic [63:0] GRF36_26_buffer [0:1];
  logic [63:0] GRF36_27_buffer [0:1];
  logic [63:0] GRF36_28_buffer [0:1];
  logic [63:0] GRF36_29_buffer [0:1];
  logic [63:0] GRF36_30_buffer [0:1];
  logic [63:0] GRF36_31_buffer [0:1];
  logic [63:0] GRF37_0_buffer [0:1];
  logic [63:0] GRF37_1_buffer [0:1];
  logic [63:0] GRF37_2_buffer [0:1];
  logic [63:0] GRF37_3_buffer [0:1];
  logic [63:0] GRF37_4_buffer [0:1];
  logic [63:0] GRF37_5_buffer [0:1];
  logic [63:0] GRF37_6_buffer [0:1];
  logic [63:0] GRF37_7_buffer [0:1];
  logic [63:0] GRF37_8_buffer [0:1];
  logic [63:0] GRF37_9_buffer [0:1];
  logic [63:0] GRF37_10_buffer [0:1];
  logic [63:0] GRF37_11_buffer [0:1];
  logic [63:0] GRF37_12_buffer [0:1];
  logic [63:0] GRF37_13_buffer [0:1];
  logic [63:0] GRF37_14_buffer [0:1];
  logic [63:0] GRF37_15_buffer [0:1];
  logic [63:0] GRF37_16_buffer [0:1];
  logic [63:0] GRF37_17_buffer [0:1];
  logic [63:0] GRF37_18_buffer [0:1];
  logic [63:0] GRF37_19_buffer [0:1];
  logic [63:0] GRF37_20_buffer [0:1];
  logic [63:0] GRF37_21_buffer [0:1];
  logic [63:0] GRF37_22_buffer [0:1];
  logic [63:0] GRF37_23_buffer [0:1];
  logic [63:0] GRF37_24_buffer [0:1];
  logic [63:0] GRF37_25_buffer [0:1];
  logic [63:0] GRF37_26_buffer [0:1];
  logic [63:0] GRF37_27_buffer [0:1];
  logic [63:0] GRF37_28_buffer [0:1];
  logic [63:0] GRF37_29_buffer [0:1];
  logic [63:0] GRF37_30_buffer [0:1];
  logic [63:0] GRF37_31_buffer [0:1];
  logic [63:0] GRF38_0_buffer [0:1];
  logic [63:0] GRF38_1_buffer [0:1];
  logic [63:0] GRF38_2_buffer [0:1];
  logic [63:0] GRF38_3_buffer [0:1];
  logic [63:0] GRF38_4_buffer [0:1];
  logic [63:0] GRF38_5_buffer [0:1];
  logic [63:0] GRF38_6_buffer [0:1];
  logic [63:0] GRF38_7_buffer [0:1];
  logic [63:0] GRF38_8_buffer [0:1];
  logic [63:0] GRF38_9_buffer [0:1];
  logic [63:0] GRF38_10_buffer [0:1];
  logic [63:0] GRF38_11_buffer [0:1];
  logic [63:0] GRF38_12_buffer [0:1];
  logic [63:0] GRF38_13_buffer [0:1];
  logic [63:0] GRF38_14_buffer [0:1];
  logic [63:0] GRF38_15_buffer [0:1];
  logic [63:0] GRF38_16_buffer [0:1];
  logic [63:0] GRF38_17_buffer [0:1];
  logic [63:0] GRF38_18_buffer [0:1];
  logic [63:0] GRF38_19_buffer [0:1];
  logic [63:0] GRF38_20_buffer [0:1];
  logic [63:0] GRF38_21_buffer [0:1];
  logic [63:0] GRF38_22_buffer [0:1];
  logic [63:0] GRF38_23_buffer [0:1];
  logic [63:0] GRF38_24_buffer [0:1];
  logic [63:0] GRF38_25_buffer [0:1];
  logic [63:0] GRF38_26_buffer [0:1];
  logic [63:0] GRF38_27_buffer [0:1];
  logic [63:0] GRF38_28_buffer [0:1];
  logic [63:0] GRF38_29_buffer [0:1];
  logic [63:0] GRF38_30_buffer [0:1];
  logic [63:0] GRF38_31_buffer [0:1];
  logic [63:0] GRF39_0_buffer [0:1];
  logic [63:0] GRF39_1_buffer [0:1];
  logic [63:0] GRF39_2_buffer [0:1];
  logic [63:0] GRF39_3_buffer [0:1];
  logic [63:0] GRF39_4_buffer [0:1];
  logic [63:0] GRF39_5_buffer [0:1];
  logic [63:0] GRF39_6_buffer [0:1];
  logic [63:0] GRF39_7_buffer [0:1];
  logic [63:0] GRF39_8_buffer [0:1];
  logic [63:0] GRF39_9_buffer [0:1];
  logic [63:0] GRF39_10_buffer [0:1];
  logic [63:0] GRF39_11_buffer [0:1];
  logic [63:0] GRF39_12_buffer [0:1];
  logic [63:0] GRF39_13_buffer [0:1];
  logic [63:0] GRF39_14_buffer [0:1];
  logic [63:0] GRF39_15_buffer [0:1];
  logic [63:0] GRF39_16_buffer [0:1];
  logic [63:0] GRF39_17_buffer [0:1];
  logic [63:0] GRF39_18_buffer [0:1];
  logic [63:0] GRF39_19_buffer [0:1];
  logic [63:0] GRF39_20_buffer [0:1];
  logic [63:0] GRF39_21_buffer [0:1];
  logic [63:0] GRF39_22_buffer [0:1];
  logic [63:0] GRF39_23_buffer [0:1];
  logic [63:0] GRF39_24_buffer [0:1];
  logic [63:0] GRF39_25_buffer [0:1];
  logic [63:0] GRF39_26_buffer [0:1];
  logic [63:0] GRF39_27_buffer [0:1];
  logic [63:0] GRF39_28_buffer [0:1];
  logic [63:0] GRF39_29_buffer [0:1];
  logic [63:0] GRF39_30_buffer [0:1];
  logic [63:0] GRF39_31_buffer [0:1];
  logic [63:0] GRF40_0_buffer [0:1];
  logic [63:0] GRF40_1_buffer [0:1];
  logic [63:0] GRF40_2_buffer [0:1];
  logic [63:0] GRF40_3_buffer [0:1];
  logic [63:0] GRF40_4_buffer [0:1];
  logic [63:0] GRF40_5_buffer [0:1];
  logic [63:0] GRF40_6_buffer [0:1];
  logic [63:0] GRF40_7_buffer [0:1];
  logic [63:0] GRF40_8_buffer [0:1];
  logic [63:0] GRF40_9_buffer [0:1];
  logic [63:0] GRF40_10_buffer [0:1];
  logic [63:0] GRF40_11_buffer [0:1];
  logic [63:0] GRF40_12_buffer [0:1];
  logic [63:0] GRF40_13_buffer [0:1];
  logic [63:0] GRF40_14_buffer [0:1];
  logic [63:0] GRF40_15_buffer [0:1];
  logic [63:0] GRF40_16_buffer [0:1];
  logic [63:0] GRF40_17_buffer [0:1];
  logic [63:0] GRF40_18_buffer [0:1];
  logic [63:0] GRF40_19_buffer [0:1];
  logic [63:0] GRF40_20_buffer [0:1];
  logic [63:0] GRF40_21_buffer [0:1];
  logic [63:0] GRF40_22_buffer [0:1];
  logic [63:0] GRF40_23_buffer [0:1];
  logic [63:0] GRF40_24_buffer [0:1];
  logic [63:0] GRF40_25_buffer [0:1];
  logic [63:0] GRF40_26_buffer [0:1];
  logic [63:0] GRF40_27_buffer [0:1];
  logic [63:0] GRF40_28_buffer [0:1];
  logic [63:0] GRF40_29_buffer [0:1];
  logic [63:0] GRF40_30_buffer [0:1];
  logic [63:0] GRF40_31_buffer [0:1];
  logic [63:0] GRF41_0_buffer [0:1];
  logic [63:0] GRF41_1_buffer [0:1];
  logic [63:0] GRF41_2_buffer [0:1];
  logic [63:0] GRF41_3_buffer [0:1];
  logic [63:0] GRF41_4_buffer [0:1];
  logic [63:0] GRF41_5_buffer [0:1];
  logic [63:0] GRF41_6_buffer [0:1];
  logic [63:0] GRF41_7_buffer [0:1];
  logic [63:0] GRF41_8_buffer [0:1];
  logic [63:0] GRF41_9_buffer [0:1];
  logic [63:0] GRF41_10_buffer [0:1];
  logic [63:0] GRF41_11_buffer [0:1];
  logic [63:0] GRF41_12_buffer [0:1];
  logic [63:0] GRF41_13_buffer [0:1];
  logic [63:0] GRF41_14_buffer [0:1];
  logic [63:0] GRF41_15_buffer [0:1];
  logic [63:0] GRF41_16_buffer [0:1];
  logic [63:0] GRF41_17_buffer [0:1];
  logic [63:0] GRF41_18_buffer [0:1];
  logic [63:0] GRF41_19_buffer [0:1];
  logic [63:0] GRF41_20_buffer [0:1];
  logic [63:0] GRF41_21_buffer [0:1];
  logic [63:0] GRF41_22_buffer [0:1];
  logic [63:0] GRF41_23_buffer [0:1];
  logic [63:0] GRF41_24_buffer [0:1];
  logic [63:0] GRF41_25_buffer [0:1];
  logic [63:0] GRF41_26_buffer [0:1];
  logic [63:0] GRF41_27_buffer [0:1];
  logic [63:0] GRF41_28_buffer [0:1];
  logic [63:0] GRF41_29_buffer [0:1];
  logic [63:0] GRF41_30_buffer [0:1];
  logic [63:0] GRF41_31_buffer [0:1];
  logic [63:0] GRF42_0_buffer [0:1];
  logic [63:0] GRF42_1_buffer [0:1];
  logic [63:0] GRF42_2_buffer [0:1];
  logic [63:0] GRF42_3_buffer [0:1];
  logic [63:0] GRF42_4_buffer [0:1];
  logic [63:0] GRF42_5_buffer [0:1];
  logic [63:0] GRF42_6_buffer [0:1];
  logic [63:0] GRF42_7_buffer [0:1];
  logic [63:0] GRF42_8_buffer [0:1];
  logic [63:0] GRF42_9_buffer [0:1];
  logic [63:0] GRF42_10_buffer [0:1];
  logic [63:0] GRF42_11_buffer [0:1];
  logic [63:0] GRF42_12_buffer [0:1];
  logic [63:0] GRF42_13_buffer [0:1];
  logic [63:0] GRF42_14_buffer [0:1];
  logic [63:0] GRF42_15_buffer [0:1];
  logic [63:0] GRF42_16_buffer [0:1];
  logic [63:0] GRF42_17_buffer [0:1];
  logic [63:0] GRF42_18_buffer [0:1];
  logic [63:0] GRF42_19_buffer [0:1];
  logic [63:0] GRF42_20_buffer [0:1];
  logic [63:0] GRF42_21_buffer [0:1];
  logic [63:0] GRF42_22_buffer [0:1];
  logic [63:0] GRF42_23_buffer [0:1];
  logic [63:0] GRF42_24_buffer [0:1];
  logic [63:0] GRF42_25_buffer [0:1];
  logic [63:0] GRF42_26_buffer [0:1];
  logic [63:0] GRF42_27_buffer [0:1];
  logic [63:0] GRF42_28_buffer [0:1];
  logic [63:0] GRF42_29_buffer [0:1];
  logic [63:0] GRF42_30_buffer [0:1];
  logic [63:0] GRF42_31_buffer [0:1];
  logic [63:0] GRF43_0_buffer [0:1];
  logic [63:0] GRF43_1_buffer [0:1];
  logic [63:0] GRF43_2_buffer [0:1];
  logic [63:0] GRF43_3_buffer [0:1];
  logic [63:0] GRF43_4_buffer [0:1];
  logic [63:0] GRF43_5_buffer [0:1];
  logic [63:0] GRF43_6_buffer [0:1];
  logic [63:0] GRF43_7_buffer [0:1];
  logic [63:0] GRF43_8_buffer [0:1];
  logic [63:0] GRF43_9_buffer [0:1];
  logic [63:0] GRF43_10_buffer [0:1];
  logic [63:0] GRF43_11_buffer [0:1];
  logic [63:0] GRF43_12_buffer [0:1];
  logic [63:0] GRF43_13_buffer [0:1];
  logic [63:0] GRF43_14_buffer [0:1];
  logic [63:0] GRF43_15_buffer [0:1];
  logic [63:0] GRF43_16_buffer [0:1];
  logic [63:0] GRF43_17_buffer [0:1];
  logic [63:0] GRF43_18_buffer [0:1];
  logic [63:0] GRF43_19_buffer [0:1];
  logic [63:0] GRF43_20_buffer [0:1];
  logic [63:0] GRF43_21_buffer [0:1];
  logic [63:0] GRF43_22_buffer [0:1];
  logic [63:0] GRF43_23_buffer [0:1];
  logic [63:0] GRF43_24_buffer [0:1];
  logic [63:0] GRF43_25_buffer [0:1];
  logic [63:0] GRF43_26_buffer [0:1];
  logic [63:0] GRF43_27_buffer [0:1];
  logic [63:0] GRF43_28_buffer [0:1];
  logic [63:0] GRF43_29_buffer [0:1];
  logic [63:0] GRF43_30_buffer [0:1];
  logic [63:0] GRF43_31_buffer [0:1];
  logic [63:0] GRF44_0_buffer [0:1];
  logic [63:0] GRF44_1_buffer [0:1];
  logic [63:0] GRF44_2_buffer [0:1];
  logic [63:0] GRF44_3_buffer [0:1];
  logic [63:0] GRF44_4_buffer [0:1];
  logic [63:0] GRF44_5_buffer [0:1];
  logic [63:0] GRF44_6_buffer [0:1];
  logic [63:0] GRF44_7_buffer [0:1];
  logic [63:0] GRF44_8_buffer [0:1];
  logic [63:0] GRF44_9_buffer [0:1];
  logic [63:0] GRF44_10_buffer [0:1];
  logic [63:0] GRF44_11_buffer [0:1];
  logic [63:0] GRF44_12_buffer [0:1];
  logic [63:0] GRF44_13_buffer [0:1];
  logic [63:0] GRF44_14_buffer [0:1];
  logic [63:0] GRF44_15_buffer [0:1];
  logic [63:0] GRF44_16_buffer [0:1];
  logic [63:0] GRF44_17_buffer [0:1];
  logic [63:0] GRF44_18_buffer [0:1];
  logic [63:0] GRF44_19_buffer [0:1];
  logic [63:0] GRF44_20_buffer [0:1];
  logic [63:0] GRF44_21_buffer [0:1];
  logic [63:0] GRF44_22_buffer [0:1];
  logic [63:0] GRF44_23_buffer [0:1];
  logic [63:0] GRF44_24_buffer [0:1];
  logic [63:0] GRF44_25_buffer [0:1];
  logic [63:0] GRF44_26_buffer [0:1];
  logic [63:0] GRF44_27_buffer [0:1];
  logic [63:0] GRF44_28_buffer [0:1];
  logic [63:0] GRF44_29_buffer [0:1];
  logic [63:0] GRF44_30_buffer [0:1];
  logic [63:0] GRF44_31_buffer [0:1];
  logic [63:0] GRF45_0_buffer [0:1];
  logic [63:0] GRF45_1_buffer [0:1];
  logic [63:0] GRF45_2_buffer [0:1];
  logic [63:0] GRF45_3_buffer [0:1];
  logic [63:0] GRF45_4_buffer [0:1];
  logic [63:0] GRF45_5_buffer [0:1];
  logic [63:0] GRF45_6_buffer [0:1];
  logic [63:0] GRF45_7_buffer [0:1];
  logic [63:0] GRF45_8_buffer [0:1];
  logic [63:0] GRF45_9_buffer [0:1];
  logic [63:0] GRF45_10_buffer [0:1];
  logic [63:0] GRF45_11_buffer [0:1];
  logic [63:0] GRF45_12_buffer [0:1];
  logic [63:0] GRF45_13_buffer [0:1];
  logic [63:0] GRF45_14_buffer [0:1];
  logic [63:0] GRF45_15_buffer [0:1];
  logic [63:0] GRF45_16_buffer [0:1];
  logic [63:0] GRF45_17_buffer [0:1];
  logic [63:0] GRF45_18_buffer [0:1];
  logic [63:0] GRF45_19_buffer [0:1];
  logic [63:0] GRF45_20_buffer [0:1];
  logic [63:0] GRF45_21_buffer [0:1];
  logic [63:0] GRF45_22_buffer [0:1];
  logic [63:0] GRF45_23_buffer [0:1];
  logic [63:0] GRF45_24_buffer [0:1];
  logic [63:0] GRF45_25_buffer [0:1];
  logic [63:0] GRF45_26_buffer [0:1];
  logic [63:0] GRF45_27_buffer [0:1];
  logic [63:0] GRF45_28_buffer [0:1];
  logic [63:0] GRF45_29_buffer [0:1];
  logic [63:0] GRF45_30_buffer [0:1];
  logic [63:0] GRF45_31_buffer [0:1];
  logic [63:0] GRF46_0_buffer [0:1];
  logic [63:0] GRF46_1_buffer [0:1];
  logic [63:0] GRF46_2_buffer [0:1];
  logic [63:0] GRF46_3_buffer [0:1];
  logic [63:0] GRF46_4_buffer [0:1];
  logic [63:0] GRF46_5_buffer [0:1];
  logic [63:0] GRF46_6_buffer [0:1];
  logic [63:0] GRF46_7_buffer [0:1];
  logic [63:0] GRF46_8_buffer [0:1];
  logic [63:0] GRF46_9_buffer [0:1];
  logic [63:0] GRF46_10_buffer [0:1];
  logic [63:0] GRF46_11_buffer [0:1];
  logic [63:0] GRF46_12_buffer [0:1];
  logic [63:0] GRF46_13_buffer [0:1];
  logic [63:0] GRF46_14_buffer [0:1];
  logic [63:0] GRF46_15_buffer [0:1];
  logic [63:0] GRF46_16_buffer [0:1];
  logic [63:0] GRF46_17_buffer [0:1];
  logic [63:0] GRF46_18_buffer [0:1];
  logic [63:0] GRF46_19_buffer [0:1];
  logic [63:0] GRF46_20_buffer [0:1];
  logic [63:0] GRF46_21_buffer [0:1];
  logic [63:0] GRF46_22_buffer [0:1];
  logic [63:0] GRF46_23_buffer [0:1];
  logic [63:0] GRF46_24_buffer [0:1];
  logic [63:0] GRF46_25_buffer [0:1];
  logic [63:0] GRF46_26_buffer [0:1];
  logic [63:0] GRF46_27_buffer [0:1];
  logic [63:0] GRF46_28_buffer [0:1];
  logic [63:0] GRF46_29_buffer [0:1];
  logic [63:0] GRF46_30_buffer [0:1];
  logic [63:0] GRF46_31_buffer [0:1];
  logic [63:0] GRF47_0_buffer [0:1];
  logic [63:0] GRF47_1_buffer [0:1];
  logic [63:0] GRF47_2_buffer [0:1];
  logic [63:0] GRF47_3_buffer [0:1];
  logic [63:0] GRF47_4_buffer [0:1];
  logic [63:0] GRF47_5_buffer [0:1];
  logic [63:0] GRF47_6_buffer [0:1];
  logic [63:0] GRF47_7_buffer [0:1];
  logic [63:0] GRF47_8_buffer [0:1];
  logic [63:0] GRF47_9_buffer [0:1];
  logic [63:0] GRF47_10_buffer [0:1];
  logic [63:0] GRF47_11_buffer [0:1];
  logic [63:0] GRF47_12_buffer [0:1];
  logic [63:0] GRF47_13_buffer [0:1];
  logic [63:0] GRF47_14_buffer [0:1];
  logic [63:0] GRF47_15_buffer [0:1];
  logic [63:0] GRF47_16_buffer [0:1];
  logic [63:0] GRF47_17_buffer [0:1];
  logic [63:0] GRF47_18_buffer [0:1];
  logic [63:0] GRF47_19_buffer [0:1];
  logic [63:0] GRF47_20_buffer [0:1];
  logic [63:0] GRF47_21_buffer [0:1];
  logic [63:0] GRF47_22_buffer [0:1];
  logic [63:0] GRF47_23_buffer [0:1];
  logic [63:0] GRF47_24_buffer [0:1];
  logic [63:0] GRF47_25_buffer [0:1];
  logic [63:0] GRF47_26_buffer [0:1];
  logic [63:0] GRF47_27_buffer [0:1];
  logic [63:0] GRF47_28_buffer [0:1];
  logic [63:0] GRF47_29_buffer [0:1];
  logic [63:0] GRF47_30_buffer [0:1];
  logic [63:0] GRF47_31_buffer [0:1];
  logic [63:0] GRF48_0_buffer [0:1];
  logic [63:0] GRF48_1_buffer [0:1];
  logic [63:0] GRF48_2_buffer [0:1];
  logic [63:0] GRF48_3_buffer [0:1];
  logic [63:0] GRF48_4_buffer [0:1];
  logic [63:0] GRF48_5_buffer [0:1];
  logic [63:0] GRF48_6_buffer [0:1];
  logic [63:0] GRF48_7_buffer [0:1];
  logic [63:0] GRF48_8_buffer [0:1];
  logic [63:0] GRF48_9_buffer [0:1];
  logic [63:0] GRF48_10_buffer [0:1];
  logic [63:0] GRF48_11_buffer [0:1];
  logic [63:0] GRF48_12_buffer [0:1];
  logic [63:0] GRF48_13_buffer [0:1];
  logic [63:0] GRF48_14_buffer [0:1];
  logic [63:0] GRF48_15_buffer [0:1];
  logic [63:0] GRF48_16_buffer [0:1];
  logic [63:0] GRF48_17_buffer [0:1];
  logic [63:0] GRF48_18_buffer [0:1];
  logic [63:0] GRF48_19_buffer [0:1];
  logic [63:0] GRF48_20_buffer [0:1];
  logic [63:0] GRF48_21_buffer [0:1];
  logic [63:0] GRF48_22_buffer [0:1];
  logic [63:0] GRF48_23_buffer [0:1];
  logic [63:0] GRF48_24_buffer [0:1];
  logic [63:0] GRF48_25_buffer [0:1];
  logic [63:0] GRF48_26_buffer [0:1];
  logic [63:0] GRF48_27_buffer [0:1];
  logic [63:0] GRF48_28_buffer [0:1];
  logic [63:0] GRF48_29_buffer [0:1];
  logic [63:0] GRF48_30_buffer [0:1];
  logic [63:0] GRF48_31_buffer [0:1];
  logic [63:0] GRF49_0_buffer [0:1];
  logic [63:0] GRF49_1_buffer [0:1];
  logic [63:0] GRF49_2_buffer [0:1];
  logic [63:0] GRF49_3_buffer [0:1];
  logic [63:0] GRF49_4_buffer [0:1];
  logic [63:0] GRF49_5_buffer [0:1];
  logic [63:0] GRF49_6_buffer [0:1];
  logic [63:0] GRF49_7_buffer [0:1];
  logic [63:0] GRF49_8_buffer [0:1];
  logic [63:0] GRF49_9_buffer [0:1];
  logic [63:0] GRF49_10_buffer [0:1];
  logic [63:0] GRF49_11_buffer [0:1];
  logic [63:0] GRF49_12_buffer [0:1];
  logic [63:0] GRF49_13_buffer [0:1];
  logic [63:0] GRF49_14_buffer [0:1];
  logic [63:0] GRF49_15_buffer [0:1];
  logic [63:0] GRF49_16_buffer [0:1];
  logic [63:0] GRF49_17_buffer [0:1];
  logic [63:0] GRF49_18_buffer [0:1];
  logic [63:0] GRF49_19_buffer [0:1];
  logic [63:0] GRF49_20_buffer [0:1];
  logic [63:0] GRF49_21_buffer [0:1];
  logic [63:0] GRF49_22_buffer [0:1];
  logic [63:0] GRF49_23_buffer [0:1];
  logic [63:0] GRF49_24_buffer [0:1];
  logic [63:0] GRF49_25_buffer [0:1];
  logic [63:0] GRF49_26_buffer [0:1];
  logic [63:0] GRF49_27_buffer [0:1];
  logic [63:0] GRF49_28_buffer [0:1];
  logic [63:0] GRF49_29_buffer [0:1];
  logic [63:0] GRF49_30_buffer [0:1];
  logic [63:0] GRF49_31_buffer [0:1];
  logic [63:0] GRF50_0_buffer [0:1];
  logic [63:0] GRF50_1_buffer [0:1];
  logic [63:0] GRF50_2_buffer [0:1];
  logic [63:0] GRF50_3_buffer [0:1];
  logic [63:0] GRF50_4_buffer [0:1];
  logic [63:0] GRF50_5_buffer [0:1];
  logic [63:0] GRF50_6_buffer [0:1];
  logic [63:0] GRF50_7_buffer [0:1];
  logic [63:0] GRF50_8_buffer [0:1];
  logic [63:0] GRF50_9_buffer [0:1];
  logic [63:0] GRF50_10_buffer [0:1];
  logic [63:0] GRF50_11_buffer [0:1];
  logic [63:0] GRF50_12_buffer [0:1];
  logic [63:0] GRF50_13_buffer [0:1];
  logic [63:0] GRF50_14_buffer [0:1];
  logic [63:0] GRF50_15_buffer [0:1];
  logic [63:0] GRF50_16_buffer [0:1];
  logic [63:0] GRF50_17_buffer [0:1];
  logic [63:0] GRF50_18_buffer [0:1];
  logic [63:0] GRF50_19_buffer [0:1];
  logic [63:0] GRF50_20_buffer [0:1];
  logic [63:0] GRF50_21_buffer [0:1];
  logic [63:0] GRF50_22_buffer [0:1];
  logic [63:0] GRF50_23_buffer [0:1];
  logic [63:0] GRF50_24_buffer [0:1];
  logic [63:0] GRF50_25_buffer [0:1];
  logic [63:0] GRF50_26_buffer [0:1];
  logic [63:0] GRF50_27_buffer [0:1];
  logic [63:0] GRF50_28_buffer [0:1];
  logic [63:0] GRF50_29_buffer [0:1];
  logic [63:0] GRF50_30_buffer [0:1];
  logic [63:0] GRF50_31_buffer [0:1];
  logic [63:0] GRF51_0_buffer [0:1];
  logic [63:0] GRF51_1_buffer [0:1];
  logic [63:0] GRF51_2_buffer [0:1];
  logic [63:0] GRF51_3_buffer [0:1];
  logic [63:0] GRF51_4_buffer [0:1];
  logic [63:0] GRF51_5_buffer [0:1];
  logic [63:0] GRF51_6_buffer [0:1];
  logic [63:0] GRF51_7_buffer [0:1];
  logic [63:0] GRF51_8_buffer [0:1];
  logic [63:0] GRF51_9_buffer [0:1];
  logic [63:0] GRF51_10_buffer [0:1];
  logic [63:0] GRF51_11_buffer [0:1];
  logic [63:0] GRF51_12_buffer [0:1];
  logic [63:0] GRF51_13_buffer [0:1];
  logic [63:0] GRF51_14_buffer [0:1];
  logic [63:0] GRF51_15_buffer [0:1];
  logic [63:0] GRF51_16_buffer [0:1];
  logic [63:0] GRF51_17_buffer [0:1];
  logic [63:0] GRF51_18_buffer [0:1];
  logic [63:0] GRF51_19_buffer [0:1];
  logic [63:0] GRF51_20_buffer [0:1];
  logic [63:0] GRF51_21_buffer [0:1];
  logic [63:0] GRF51_22_buffer [0:1];
  logic [63:0] GRF51_23_buffer [0:1];
  logic [63:0] GRF51_24_buffer [0:1];
  logic [63:0] GRF51_25_buffer [0:1];
  logic [63:0] GRF51_26_buffer [0:1];
  logic [63:0] GRF51_27_buffer [0:1];
  logic [63:0] GRF51_28_buffer [0:1];
  logic [63:0] GRF51_29_buffer [0:1];
  logic [63:0] GRF51_30_buffer [0:1];
  logic [63:0] GRF51_31_buffer [0:1];
  logic [63:0] GRF52_0_buffer [0:1];
  logic [63:0] GRF52_1_buffer [0:1];
  logic [63:0] GRF52_2_buffer [0:1];
  logic [63:0] GRF52_3_buffer [0:1];
  logic [63:0] GRF52_4_buffer [0:1];
  logic [63:0] GRF52_5_buffer [0:1];
  logic [63:0] GRF52_6_buffer [0:1];
  logic [63:0] GRF52_7_buffer [0:1];
  logic [63:0] GRF52_8_buffer [0:1];
  logic [63:0] GRF52_9_buffer [0:1];
  logic [63:0] GRF52_10_buffer [0:1];
  logic [63:0] GRF52_11_buffer [0:1];
  logic [63:0] GRF52_12_buffer [0:1];
  logic [63:0] GRF52_13_buffer [0:1];
  logic [63:0] GRF52_14_buffer [0:1];
  logic [63:0] GRF52_15_buffer [0:1];
  logic [63:0] GRF52_16_buffer [0:1];
  logic [63:0] GRF52_17_buffer [0:1];
  logic [63:0] GRF52_18_buffer [0:1];
  logic [63:0] GRF52_19_buffer [0:1];
  logic [63:0] GRF52_20_buffer [0:1];
  logic [63:0] GRF52_21_buffer [0:1];
  logic [63:0] GRF52_22_buffer [0:1];
  logic [63:0] GRF52_23_buffer [0:1];
  logic [63:0] GRF52_24_buffer [0:1];
  logic [63:0] GRF52_25_buffer [0:1];
  logic [63:0] GRF52_26_buffer [0:1];
  logic [63:0] GRF52_27_buffer [0:1];
  logic [63:0] GRF52_28_buffer [0:1];
  logic [63:0] GRF52_29_buffer [0:1];
  logic [63:0] GRF52_30_buffer [0:1];
  logic [63:0] GRF52_31_buffer [0:1];
  logic [63:0] GRF53_0_buffer [0:1];
  logic [63:0] GRF53_1_buffer [0:1];
  logic [63:0] GRF53_2_buffer [0:1];
  logic [63:0] GRF53_3_buffer [0:1];
  logic [63:0] GRF53_4_buffer [0:1];
  logic [63:0] GRF53_5_buffer [0:1];
  logic [63:0] GRF53_6_buffer [0:1];
  logic [63:0] GRF53_7_buffer [0:1];
  logic [63:0] GRF53_8_buffer [0:1];
  logic [63:0] GRF53_9_buffer [0:1];
  logic [63:0] GRF53_10_buffer [0:1];
  logic [63:0] GRF53_11_buffer [0:1];
  logic [63:0] GRF53_12_buffer [0:1];
  logic [63:0] GRF53_13_buffer [0:1];
  logic [63:0] GRF53_14_buffer [0:1];
  logic [63:0] GRF53_15_buffer [0:1];
  logic [63:0] GRF53_16_buffer [0:1];
  logic [63:0] GRF53_17_buffer [0:1];
  logic [63:0] GRF53_18_buffer [0:1];
  logic [63:0] GRF53_19_buffer [0:1];
  logic [63:0] GRF53_20_buffer [0:1];
  logic [63:0] GRF53_21_buffer [0:1];
  logic [63:0] GRF53_22_buffer [0:1];
  logic [63:0] GRF53_23_buffer [0:1];
  logic [63:0] GRF53_24_buffer [0:1];
  logic [63:0] GRF53_25_buffer [0:1];
  logic [63:0] GRF53_26_buffer [0:1];
  logic [63:0] GRF53_27_buffer [0:1];
  logic [63:0] GRF53_28_buffer [0:1];
  logic [63:0] GRF53_29_buffer [0:1];
  logic [63:0] GRF53_30_buffer [0:1];
  logic [63:0] GRF53_31_buffer [0:1];
  logic [63:0] GRF54_0_buffer [0:1];
  logic [63:0] GRF54_1_buffer [0:1];
  logic [63:0] GRF54_2_buffer [0:1];
  logic [63:0] GRF54_3_buffer [0:1];
  logic [63:0] GRF54_4_buffer [0:1];
  logic [63:0] GRF54_5_buffer [0:1];
  logic [63:0] GRF54_6_buffer [0:1];
  logic [63:0] GRF54_7_buffer [0:1];
  logic [63:0] GRF54_8_buffer [0:1];
  logic [63:0] GRF54_9_buffer [0:1];
  logic [63:0] GRF54_10_buffer [0:1];
  logic [63:0] GRF54_11_buffer [0:1];
  logic [63:0] GRF54_12_buffer [0:1];
  logic [63:0] GRF54_13_buffer [0:1];
  logic [63:0] GRF54_14_buffer [0:1];
  logic [63:0] GRF54_15_buffer [0:1];
  logic [63:0] GRF54_16_buffer [0:1];
  logic [63:0] GRF54_17_buffer [0:1];
  logic [63:0] GRF54_18_buffer [0:1];
  logic [63:0] GRF54_19_buffer [0:1];
  logic [63:0] GRF54_20_buffer [0:1];
  logic [63:0] GRF54_21_buffer [0:1];
  logic [63:0] GRF54_22_buffer [0:1];
  logic [63:0] GRF54_23_buffer [0:1];
  logic [63:0] GRF54_24_buffer [0:1];
  logic [63:0] GRF54_25_buffer [0:1];
  logic [63:0] GRF54_26_buffer [0:1];
  logic [63:0] GRF54_27_buffer [0:1];
  logic [63:0] GRF54_28_buffer [0:1];
  logic [63:0] GRF54_29_buffer [0:1];
  logic [63:0] GRF54_30_buffer [0:1];
  logic [63:0] GRF54_31_buffer [0:1];
  logic [63:0] GRF55_0_buffer [0:1];
  logic [63:0] GRF55_1_buffer [0:1];
  logic [63:0] GRF55_2_buffer [0:1];
  logic [63:0] GRF55_3_buffer [0:1];
  logic [63:0] GRF55_4_buffer [0:1];
  logic [63:0] GRF55_5_buffer [0:1];
  logic [63:0] GRF55_6_buffer [0:1];
  logic [63:0] GRF55_7_buffer [0:1];
  logic [63:0] GRF55_8_buffer [0:1];
  logic [63:0] GRF55_9_buffer [0:1];
  logic [63:0] GRF55_10_buffer [0:1];
  logic [63:0] GRF55_11_buffer [0:1];
  logic [63:0] GRF55_12_buffer [0:1];
  logic [63:0] GRF55_13_buffer [0:1];
  logic [63:0] GRF55_14_buffer [0:1];
  logic [63:0] GRF55_15_buffer [0:1];
  logic [63:0] GRF55_16_buffer [0:1];
  logic [63:0] GRF55_17_buffer [0:1];
  logic [63:0] GRF55_18_buffer [0:1];
  logic [63:0] GRF55_19_buffer [0:1];
  logic [63:0] GRF55_20_buffer [0:1];
  logic [63:0] GRF55_21_buffer [0:1];
  logic [63:0] GRF55_22_buffer [0:1];
  logic [63:0] GRF55_23_buffer [0:1];
  logic [63:0] GRF55_24_buffer [0:1];
  logic [63:0] GRF55_25_buffer [0:1];
  logic [63:0] GRF55_26_buffer [0:1];
  logic [63:0] GRF55_27_buffer [0:1];
  logic [63:0] GRF55_28_buffer [0:1];
  logic [63:0] GRF55_29_buffer [0:1];
  logic [63:0] GRF55_30_buffer [0:1];
  logic [63:0] GRF55_31_buffer [0:1];
  logic [63:0] GRF56_0_buffer [0:1];
  logic [63:0] GRF56_1_buffer [0:1];
  logic [63:0] GRF56_2_buffer [0:1];
  logic [63:0] GRF56_3_buffer [0:1];
  logic [63:0] GRF56_4_buffer [0:1];
  logic [63:0] GRF56_5_buffer [0:1];
  logic [63:0] GRF56_6_buffer [0:1];
  logic [63:0] GRF56_7_buffer [0:1];
  logic [63:0] GRF56_8_buffer [0:1];
  logic [63:0] GRF56_9_buffer [0:1];
  logic [63:0] GRF56_10_buffer [0:1];
  logic [63:0] GRF56_11_buffer [0:1];
  logic [63:0] GRF56_12_buffer [0:1];
  logic [63:0] GRF56_13_buffer [0:1];
  logic [63:0] GRF56_14_buffer [0:1];
  logic [63:0] GRF56_15_buffer [0:1];
  logic [63:0] GRF56_16_buffer [0:1];
  logic [63:0] GRF56_17_buffer [0:1];
  logic [63:0] GRF56_18_buffer [0:1];
  logic [63:0] GRF56_19_buffer [0:1];
  logic [63:0] GRF56_20_buffer [0:1];
  logic [63:0] GRF56_21_buffer [0:1];
  logic [63:0] GRF56_22_buffer [0:1];
  logic [63:0] GRF56_23_buffer [0:1];
  logic [63:0] GRF56_24_buffer [0:1];
  logic [63:0] GRF56_25_buffer [0:1];
  logic [63:0] GRF56_26_buffer [0:1];
  logic [63:0] GRF56_27_buffer [0:1];
  logic [63:0] GRF56_28_buffer [0:1];
  logic [63:0] GRF56_29_buffer [0:1];
  logic [63:0] GRF56_30_buffer [0:1];
  logic [63:0] GRF56_31_buffer [0:1];
  logic [63:0] GRF57_0_buffer [0:1];
  logic [63:0] GRF57_1_buffer [0:1];
  logic [63:0] GRF57_2_buffer [0:1];
  logic [63:0] GRF57_3_buffer [0:1];
  logic [63:0] GRF57_4_buffer [0:1];
  logic [63:0] GRF57_5_buffer [0:1];
  logic [63:0] GRF57_6_buffer [0:1];
  logic [63:0] GRF57_7_buffer [0:1];
  logic [63:0] GRF57_8_buffer [0:1];
  logic [63:0] GRF57_9_buffer [0:1];
  logic [63:0] GRF57_10_buffer [0:1];
  logic [63:0] GRF57_11_buffer [0:1];
  logic [63:0] GRF57_12_buffer [0:1];
  logic [63:0] GRF57_13_buffer [0:1];
  logic [63:0] GRF57_14_buffer [0:1];
  logic [63:0] GRF57_15_buffer [0:1];
  logic [63:0] GRF57_16_buffer [0:1];
  logic [63:0] GRF57_17_buffer [0:1];
  logic [63:0] GRF57_18_buffer [0:1];
  logic [63:0] GRF57_19_buffer [0:1];
  logic [63:0] GRF57_20_buffer [0:1];
  logic [63:0] GRF57_21_buffer [0:1];
  logic [63:0] GRF57_22_buffer [0:1];
  logic [63:0] GRF57_23_buffer [0:1];
  logic [63:0] GRF57_24_buffer [0:1];
  logic [63:0] GRF57_25_buffer [0:1];
  logic [63:0] GRF57_26_buffer [0:1];
  logic [63:0] GRF57_27_buffer [0:1];
  logic [63:0] GRF57_28_buffer [0:1];
  logic [63:0] GRF57_29_buffer [0:1];
  logic [63:0] GRF57_30_buffer [0:1];
  logic [63:0] GRF57_31_buffer [0:1];
  logic [63:0] GRF58_0_buffer [0:1];
  logic [63:0] GRF58_1_buffer [0:1];
  logic [63:0] GRF58_2_buffer [0:1];
  logic [63:0] GRF58_3_buffer [0:1];
  logic [63:0] GRF58_4_buffer [0:1];
  logic [63:0] GRF58_5_buffer [0:1];
  logic [63:0] GRF58_6_buffer [0:1];
  logic [63:0] GRF58_7_buffer [0:1];
  logic [63:0] GRF58_8_buffer [0:1];
  logic [63:0] GRF58_9_buffer [0:1];
  logic [63:0] GRF58_10_buffer [0:1];
  logic [63:0] GRF58_11_buffer [0:1];
  logic [63:0] GRF58_12_buffer [0:1];
  logic [63:0] GRF58_13_buffer [0:1];
  logic [63:0] GRF58_14_buffer [0:1];
  logic [63:0] GRF58_15_buffer [0:1];
  logic [63:0] GRF58_16_buffer [0:1];
  logic [63:0] GRF58_17_buffer [0:1];
  logic [63:0] GRF58_18_buffer [0:1];
  logic [63:0] GRF58_19_buffer [0:1];
  logic [63:0] GRF58_20_buffer [0:1];
  logic [63:0] GRF58_21_buffer [0:1];
  logic [63:0] GRF58_22_buffer [0:1];
  logic [63:0] GRF58_23_buffer [0:1];
  logic [63:0] GRF58_24_buffer [0:1];
  logic [63:0] GRF58_25_buffer [0:1];
  logic [63:0] GRF58_26_buffer [0:1];
  logic [63:0] GRF58_27_buffer [0:1];
  logic [63:0] GRF58_28_buffer [0:1];
  logic [63:0] GRF58_29_buffer [0:1];
  logic [63:0] GRF58_30_buffer [0:1];
  logic [63:0] GRF58_31_buffer [0:1];
  logic [63:0] GRF59_0_buffer [0:1];
  logic [63:0] GRF59_1_buffer [0:1];
  logic [63:0] GRF59_2_buffer [0:1];
  logic [63:0] GRF59_3_buffer [0:1];
  logic [63:0] GRF59_4_buffer [0:1];
  logic [63:0] GRF59_5_buffer [0:1];
  logic [63:0] GRF59_6_buffer [0:1];
  logic [63:0] GRF59_7_buffer [0:1];
  logic [63:0] GRF59_8_buffer [0:1];
  logic [63:0] GRF59_9_buffer [0:1];
  logic [63:0] GRF59_10_buffer [0:1];
  logic [63:0] GRF59_11_buffer [0:1];
  logic [63:0] GRF59_12_buffer [0:1];
  logic [63:0] GRF59_13_buffer [0:1];
  logic [63:0] GRF59_14_buffer [0:1];
  logic [63:0] GRF59_15_buffer [0:1];
  logic [63:0] GRF59_16_buffer [0:1];
  logic [63:0] GRF59_17_buffer [0:1];
  logic [63:0] GRF59_18_buffer [0:1];
  logic [63:0] GRF59_19_buffer [0:1];
  logic [63:0] GRF59_20_buffer [0:1];
  logic [63:0] GRF59_21_buffer [0:1];
  logic [63:0] GRF59_22_buffer [0:1];
  logic [63:0] GRF59_23_buffer [0:1];
  logic [63:0] GRF59_24_buffer [0:1];
  logic [63:0] GRF59_25_buffer [0:1];
  logic [63:0] GRF59_26_buffer [0:1];
  logic [63:0] GRF59_27_buffer [0:1];
  logic [63:0] GRF59_28_buffer [0:1];
  logic [63:0] GRF59_29_buffer [0:1];
  logic [63:0] GRF59_30_buffer [0:1];
  logic [63:0] GRF59_31_buffer [0:1];
  logic [63:0] GRF60_0_buffer [0:1];
  logic [63:0] GRF60_1_buffer [0:1];
  logic [63:0] GRF60_2_buffer [0:1];
  logic [63:0] GRF60_3_buffer [0:1];
  logic [63:0] GRF60_4_buffer [0:1];
  logic [63:0] GRF60_5_buffer [0:1];
  logic [63:0] GRF60_6_buffer [0:1];
  logic [63:0] GRF60_7_buffer [0:1];
  logic [63:0] GRF60_8_buffer [0:1];
  logic [63:0] GRF60_9_buffer [0:1];
  logic [63:0] GRF60_10_buffer [0:1];
  logic [63:0] GRF60_11_buffer [0:1];
  logic [63:0] GRF60_12_buffer [0:1];
  logic [63:0] GRF60_13_buffer [0:1];
  logic [63:0] GRF60_14_buffer [0:1];
  logic [63:0] GRF60_15_buffer [0:1];
  logic [63:0] GRF60_16_buffer [0:1];
  logic [63:0] GRF60_17_buffer [0:1];
  logic [63:0] GRF60_18_buffer [0:1];
  logic [63:0] GRF60_19_buffer [0:1];
  logic [63:0] GRF60_20_buffer [0:1];
  logic [63:0] GRF60_21_buffer [0:1];
  logic [63:0] GRF60_22_buffer [0:1];
  logic [63:0] GRF60_23_buffer [0:1];
  logic [63:0] GRF60_24_buffer [0:1];
  logic [63:0] GRF60_25_buffer [0:1];
  logic [63:0] GRF60_26_buffer [0:1];
  logic [63:0] GRF60_27_buffer [0:1];
  logic [63:0] GRF60_28_buffer [0:1];
  logic [63:0] GRF60_29_buffer [0:1];
  logic [63:0] GRF60_30_buffer [0:1];
  logic [63:0] GRF60_31_buffer [0:1];
  logic [63:0] GRF61_0_buffer [0:1];
  logic [63:0] GRF61_1_buffer [0:1];
  logic [63:0] GRF61_2_buffer [0:1];
  logic [63:0] GRF61_3_buffer [0:1];
  logic [63:0] GRF61_4_buffer [0:1];
  logic [63:0] GRF61_5_buffer [0:1];
  logic [63:0] GRF61_6_buffer [0:1];
  logic [63:0] GRF61_7_buffer [0:1];
  logic [63:0] GRF61_8_buffer [0:1];
  logic [63:0] GRF61_9_buffer [0:1];
  logic [63:0] GRF61_10_buffer [0:1];
  logic [63:0] GRF61_11_buffer [0:1];
  logic [63:0] GRF61_12_buffer [0:1];
  logic [63:0] GRF61_13_buffer [0:1];
  logic [63:0] GRF61_14_buffer [0:1];
  logic [63:0] GRF61_15_buffer [0:1];
  logic [63:0] GRF61_16_buffer [0:1];
  logic [63:0] GRF61_17_buffer [0:1];
  logic [63:0] GRF61_18_buffer [0:1];
  logic [63:0] GRF61_19_buffer [0:1];
  logic [63:0] GRF61_20_buffer [0:1];
  logic [63:0] GRF61_21_buffer [0:1];
  logic [63:0] GRF61_22_buffer [0:1];
  logic [63:0] GRF61_23_buffer [0:1];
  logic [63:0] GRF61_24_buffer [0:1];
  logic [63:0] GRF61_25_buffer [0:1];
  logic [63:0] GRF61_26_buffer [0:1];
  logic [63:0] GRF61_27_buffer [0:1];
  logic [63:0] GRF61_28_buffer [0:1];
  logic [63:0] GRF61_29_buffer [0:1];
  logic [63:0] GRF61_30_buffer [0:1];
  logic [63:0] GRF61_31_buffer [0:1];
  logic [63:0] GRF62_0_buffer [0:1];
  logic [63:0] GRF62_1_buffer [0:1];
  logic [63:0] GRF62_2_buffer [0:1];
  logic [63:0] GRF62_3_buffer [0:1];
  logic [63:0] GRF62_4_buffer [0:1];
  logic [63:0] GRF62_5_buffer [0:1];
  logic [63:0] GRF62_6_buffer [0:1];
  logic [63:0] GRF62_7_buffer [0:1];
  logic [63:0] GRF62_8_buffer [0:1];
  logic [63:0] GRF62_9_buffer [0:1];
  logic [63:0] GRF62_10_buffer [0:1];
  logic [63:0] GRF62_11_buffer [0:1];
  logic [63:0] GRF62_12_buffer [0:1];
  logic [63:0] GRF62_13_buffer [0:1];
  logic [63:0] GRF62_14_buffer [0:1];
  logic [63:0] GRF62_15_buffer [0:1];
  logic [63:0] GRF62_16_buffer [0:1];
  logic [63:0] GRF62_17_buffer [0:1];
  logic [63:0] GRF62_18_buffer [0:1];
  logic [63:0] GRF62_19_buffer [0:1];
  logic [63:0] GRF62_20_buffer [0:1];
  logic [63:0] GRF62_21_buffer [0:1];
  logic [63:0] GRF62_22_buffer [0:1];
  logic [63:0] GRF62_23_buffer [0:1];
  logic [63:0] GRF62_24_buffer [0:1];
  logic [63:0] GRF62_25_buffer [0:1];
  logic [63:0] GRF62_26_buffer [0:1];
  logic [63:0] GRF62_27_buffer [0:1];
  logic [63:0] GRF62_28_buffer [0:1];
  logic [63:0] GRF62_29_buffer [0:1];
  logic [63:0] GRF62_30_buffer [0:1];
  logic [63:0] GRF62_31_buffer [0:1];
  logic [63:0] GRF63_0_buffer [0:1];
  logic [63:0] GRF63_1_buffer [0:1];
  logic [63:0] GRF63_2_buffer [0:1];
  logic [63:0] GRF63_3_buffer [0:1];
  logic [63:0] GRF63_4_buffer [0:1];
  logic [63:0] GRF63_5_buffer [0:1];
  logic [63:0] GRF63_6_buffer [0:1];
  logic [63:0] GRF63_7_buffer [0:1];
  logic [63:0] GRF63_8_buffer [0:1];
  logic [63:0] GRF63_9_buffer [0:1];
  logic [63:0] GRF63_10_buffer [0:1];
  logic [63:0] GRF63_11_buffer [0:1];
  logic [63:0] GRF63_12_buffer [0:1];
  logic [63:0] GRF63_13_buffer [0:1];
  logic [63:0] GRF63_14_buffer [0:1];
  logic [63:0] GRF63_15_buffer [0:1];
  logic [63:0] GRF63_16_buffer [0:1];
  logic [63:0] GRF63_17_buffer [0:1];
  logic [63:0] GRF63_18_buffer [0:1];
  logic [63:0] GRF63_19_buffer [0:1];
  logic [63:0] GRF63_20_buffer [0:1];
  logic [63:0] GRF63_21_buffer [0:1];
  logic [63:0] GRF63_22_buffer [0:1];
  logic [63:0] GRF63_23_buffer [0:1];
  logic [63:0] GRF63_24_buffer [0:1];
  logic [63:0] GRF63_25_buffer [0:1];
  logic [63:0] GRF63_26_buffer [0:1];
  logic [63:0] GRF63_27_buffer [0:1];
  logic [63:0] GRF63_28_buffer [0:1];
  logic [63:0] GRF63_29_buffer [0:1];
  logic [63:0] GRF63_30_buffer [0:1];
  logic [63:0] GRF63_31_buffer [0:1];

  // initiate warp signals (1 if there is a change in one of the buffers)
  logic warp0_sig;
  logic warp1_sig;
  logic warp2_sig;
  logic warp3_sig;
  logic warp4_sig;
  logic warp5_sig;
  logic warp6_sig;
  logic warp7_sig;


  // Initialize the output tracker file
  initial begin
    f = $fopen("h_tracker.txt", "w");
    $fwrite(f, "=====================================================\n");
    $fwrite(f, "              Harmonica Tracker v1");
    $fwrite(f, " \n=====================================================\n\n");

  end


  // Need to differentiate between different warps time instruction and changes to memory and registers

  // Put information into the buffer // FIXME, code bloat // for loop  -- syntax for printing is not correct, so i just copied and paste from C++ code // FIXME
  always @ (edge clk) begin
    GRF0_0_buffer[clk] = GRF0[0];
    GRF0_1_buffer[clk] = GRF0[1];
    GRF0_2_buffer[clk] = GRF0[2];
    GRF0_3_buffer[clk] = GRF0[3];
    GRF0_4_buffer[clk] = GRF0[4];
    GRF0_5_buffer[clk] = GRF0[5];
    GRF0_6_buffer[clk] = GRF0[6];
    GRF0_7_buffer[clk] = GRF0[7];
    GRF0_8_buffer[clk] = GRF0[8];
    GRF0_9_buffer[clk] = GRF0[9];
    GRF0_10_buffer[clk] = GRF0[10];
    GRF0_11_buffer[clk] = GRF0[11];
    GRF0_12_buffer[clk] = GRF0[12];
    GRF0_13_buffer[clk] = GRF0[13];
    GRF0_14_buffer[clk] = GRF0[14];
    GRF0_15_buffer[clk] = GRF0[15];
    GRF0_16_buffer[clk] = GRF0[16];
    GRF0_17_buffer[clk] = GRF0[17];
    GRF0_18_buffer[clk] = GRF0[18];
    GRF0_19_buffer[clk] = GRF0[19];
    GRF0_20_buffer[clk] = GRF0[20];
    GRF0_21_buffer[clk] = GRF0[21];
    GRF0_22_buffer[clk] = GRF0[22];
    GRF0_23_buffer[clk] = GRF0[23];
    GRF0_24_buffer[clk] = GRF0[24];
    GRF0_25_buffer[clk] = GRF0[25];
    GRF0_26_buffer[clk] = GRF0[26];
    GRF0_27_buffer[clk] = GRF0[27];
    GRF0_28_buffer[clk] = GRF0[28];
    GRF0_29_buffer[clk] = GRF0[29];
    GRF0_30_buffer[clk] = GRF0[30];
    GRF0_31_buffer[clk] = GRF0[31];
    GRF1_0_buffer[clk] = GRF1[0];
    GRF1_1_buffer[clk] = GRF1[1];
    GRF1_2_buffer[clk] = GRF1[2];
    GRF1_3_buffer[clk] = GRF1[3];
    GRF1_4_buffer[clk] = GRF1[4];
    GRF1_5_buffer[clk] = GRF1[5];
    GRF1_6_buffer[clk] = GRF1[6];
    GRF1_7_buffer[clk] = GRF1[7];
    GRF1_8_buffer[clk] = GRF1[8];
    GRF1_9_buffer[clk] = GRF1[9];
    GRF1_10_buffer[clk] = GRF1[10];
    GRF1_11_buffer[clk] = GRF1[11];
    GRF1_12_buffer[clk] = GRF1[12];
    GRF1_13_buffer[clk] = GRF1[13];
    GRF1_14_buffer[clk] = GRF1[14];
    GRF1_15_buffer[clk] = GRF1[15];
    GRF1_16_buffer[clk] = GRF1[16];
    GRF1_17_buffer[clk] = GRF1[17];
    GRF1_18_buffer[clk] = GRF1[18];
    GRF1_19_buffer[clk] = GRF1[19];
    GRF1_20_buffer[clk] = GRF1[20];
    GRF1_21_buffer[clk] = GRF1[21];
    GRF1_22_buffer[clk] = GRF1[22];
    GRF1_23_buffer[clk] = GRF1[23];
    GRF1_24_buffer[clk] = GRF1[24];
    GRF1_25_buffer[clk] = GRF1[25];
    GRF1_26_buffer[clk] = GRF1[26];
    GRF1_27_buffer[clk] = GRF1[27];
    GRF1_28_buffer[clk] = GRF1[28];
    GRF1_29_buffer[clk] = GRF1[29];
    GRF1_30_buffer[clk] = GRF1[30];
    GRF1_31_buffer[clk] = GRF1[31];
    GRF2_0_buffer[clk] = GRF2[0];
    GRF2_1_buffer[clk] = GRF2[1];
    GRF2_2_buffer[clk] = GRF2[2];
    GRF2_3_buffer[clk] = GRF2[3];
    GRF2_4_buffer[clk] = GRF2[4];
    GRF2_5_buffer[clk] = GRF2[5];
    GRF2_6_buffer[clk] = GRF2[6];
    GRF2_7_buffer[clk] = GRF2[7];
    GRF2_8_buffer[clk] = GRF2[8];
    GRF2_9_buffer[clk] = GRF2[9];
    GRF2_10_buffer[clk] = GRF2[10];
    GRF2_11_buffer[clk] = GRF2[11];
    GRF2_12_buffer[clk] = GRF2[12];
    GRF2_13_buffer[clk] = GRF2[13];
    GRF2_14_buffer[clk] = GRF2[14];
    GRF2_15_buffer[clk] = GRF2[15];
    GRF2_16_buffer[clk] = GRF2[16];
    GRF2_17_buffer[clk] = GRF2[17];
    GRF2_18_buffer[clk] = GRF2[18];
    GRF2_19_buffer[clk] = GRF2[19];
    GRF2_20_buffer[clk] = GRF2[20];
    GRF2_21_buffer[clk] = GRF2[21];
    GRF2_22_buffer[clk] = GRF2[22];
    GRF2_23_buffer[clk] = GRF2[23];
    GRF2_24_buffer[clk] = GRF2[24];
    GRF2_25_buffer[clk] = GRF2[25];
    GRF2_26_buffer[clk] = GRF2[26];
    GRF2_27_buffer[clk] = GRF2[27];
    GRF2_28_buffer[clk] = GRF2[28];
    GRF2_29_buffer[clk] = GRF2[29];
    GRF2_30_buffer[clk] = GRF2[30];
    GRF2_31_buffer[clk] = GRF2[31];
    GRF3_0_buffer[clk] = GRF3[0];
    GRF3_1_buffer[clk] = GRF3[1];
    GRF3_2_buffer[clk] = GRF3[2];
    GRF3_3_buffer[clk] = GRF3[3];
    GRF3_4_buffer[clk] = GRF3[4];
    GRF3_5_buffer[clk] = GRF3[5];
    GRF3_6_buffer[clk] = GRF3[6];
    GRF3_7_buffer[clk] = GRF3[7];
    GRF3_8_buffer[clk] = GRF3[8];
    GRF3_9_buffer[clk] = GRF3[9];
    GRF3_10_buffer[clk] = GRF3[10];
    GRF3_11_buffer[clk] = GRF3[11];
    GRF3_12_buffer[clk] = GRF3[12];
    GRF3_13_buffer[clk] = GRF3[13];
    GRF3_14_buffer[clk] = GRF3[14];
    GRF3_15_buffer[clk] = GRF3[15];
    GRF3_16_buffer[clk] = GRF3[16];
    GRF3_17_buffer[clk] = GRF3[17];
    GRF3_18_buffer[clk] = GRF3[18];
    GRF3_19_buffer[clk] = GRF3[19];
    GRF3_20_buffer[clk] = GRF3[20];
    GRF3_21_buffer[clk] = GRF3[21];
    GRF3_22_buffer[clk] = GRF3[22];
    GRF3_23_buffer[clk] = GRF3[23];
    GRF3_24_buffer[clk] = GRF3[24];
    GRF3_25_buffer[clk] = GRF3[25];
    GRF3_26_buffer[clk] = GRF3[26];
    GRF3_27_buffer[clk] = GRF3[27];
    GRF3_28_buffer[clk] = GRF3[28];
    GRF3_29_buffer[clk] = GRF3[29];
    GRF3_30_buffer[clk] = GRF3[30];
    GRF3_31_buffer[clk] = GRF3[31];
    GRF4_0_buffer[clk] = GRF4[0];
    GRF4_1_buffer[clk] = GRF4[1];
    GRF4_2_buffer[clk] = GRF4[2];
    GRF4_3_buffer[clk] = GRF4[3];
    GRF4_4_buffer[clk] = GRF4[4];
    GRF4_5_buffer[clk] = GRF4[5];
    GRF4_6_buffer[clk] = GRF4[6];
    GRF4_7_buffer[clk] = GRF4[7];
    GRF4_8_buffer[clk] = GRF4[8];
    GRF4_9_buffer[clk] = GRF4[9];
    GRF4_10_buffer[clk] = GRF4[10];
    GRF4_11_buffer[clk] = GRF4[11];
    GRF4_12_buffer[clk] = GRF4[12];
    GRF4_13_buffer[clk] = GRF4[13];
    GRF4_14_buffer[clk] = GRF4[14];
    GRF4_15_buffer[clk] = GRF4[15];
    GRF4_16_buffer[clk] = GRF4[16];
    GRF4_17_buffer[clk] = GRF4[17];
    GRF4_18_buffer[clk] = GRF4[18];
    GRF4_19_buffer[clk] = GRF4[19];
    GRF4_20_buffer[clk] = GRF4[20];
    GRF4_21_buffer[clk] = GRF4[21];
    GRF4_22_buffer[clk] = GRF4[22];
    GRF4_23_buffer[clk] = GRF4[23];
    GRF4_24_buffer[clk] = GRF4[24];
    GRF4_25_buffer[clk] = GRF4[25];
    GRF4_26_buffer[clk] = GRF4[26];
    GRF4_27_buffer[clk] = GRF4[27];
    GRF4_28_buffer[clk] = GRF4[28];
    GRF4_29_buffer[clk] = GRF4[29];
    GRF4_30_buffer[clk] = GRF4[30];
    GRF4_31_buffer[clk] = GRF4[31];
    GRF5_0_buffer[clk] = GRF5[0];
    GRF5_1_buffer[clk] = GRF5[1];
    GRF5_2_buffer[clk] = GRF5[2];
    GRF5_3_buffer[clk] = GRF5[3];
    GRF5_4_buffer[clk] = GRF5[4];
    GRF5_5_buffer[clk] = GRF5[5];
    GRF5_6_buffer[clk] = GRF5[6];
    GRF5_7_buffer[clk] = GRF5[7];
    GRF5_8_buffer[clk] = GRF5[8];
    GRF5_9_buffer[clk] = GRF5[9];
    GRF5_10_buffer[clk] = GRF5[10];
    GRF5_11_buffer[clk] = GRF5[11];
    GRF5_12_buffer[clk] = GRF5[12];
    GRF5_13_buffer[clk] = GRF5[13];
    GRF5_14_buffer[clk] = GRF5[14];
    GRF5_15_buffer[clk] = GRF5[15];
    GRF5_16_buffer[clk] = GRF5[16];
    GRF5_17_buffer[clk] = GRF5[17];
    GRF5_18_buffer[clk] = GRF5[18];
    GRF5_19_buffer[clk] = GRF5[19];
    GRF5_20_buffer[clk] = GRF5[20];
    GRF5_21_buffer[clk] = GRF5[21];
    GRF5_22_buffer[clk] = GRF5[22];
    GRF5_23_buffer[clk] = GRF5[23];
    GRF5_24_buffer[clk] = GRF5[24];
    GRF5_25_buffer[clk] = GRF5[25];
    GRF5_26_buffer[clk] = GRF5[26];
    GRF5_27_buffer[clk] = GRF5[27];
    GRF5_28_buffer[clk] = GRF5[28];
    GRF5_29_buffer[clk] = GRF5[29];
    GRF5_30_buffer[clk] = GRF5[30];
    GRF5_31_buffer[clk] = GRF5[31];
    GRF6_0_buffer[clk] = GRF6[0];
    GRF6_1_buffer[clk] = GRF6[1];
    GRF6_2_buffer[clk] = GRF6[2];
    GRF6_3_buffer[clk] = GRF6[3];
    GRF6_4_buffer[clk] = GRF6[4];
    GRF6_5_buffer[clk] = GRF6[5];
    GRF6_6_buffer[clk] = GRF6[6];
    GRF6_7_buffer[clk] = GRF6[7];
    GRF6_8_buffer[clk] = GRF6[8];
    GRF6_9_buffer[clk] = GRF6[9];
    GRF6_10_buffer[clk] = GRF6[10];
    GRF6_11_buffer[clk] = GRF6[11];
    GRF6_12_buffer[clk] = GRF6[12];
    GRF6_13_buffer[clk] = GRF6[13];
    GRF6_14_buffer[clk] = GRF6[14];
    GRF6_15_buffer[clk] = GRF6[15];
    GRF6_16_buffer[clk] = GRF6[16];
    GRF6_17_buffer[clk] = GRF6[17];
    GRF6_18_buffer[clk] = GRF6[18];
    GRF6_19_buffer[clk] = GRF6[19];
    GRF6_20_buffer[clk] = GRF6[20];
    GRF6_21_buffer[clk] = GRF6[21];
    GRF6_22_buffer[clk] = GRF6[22];
    GRF6_23_buffer[clk] = GRF6[23];
    GRF6_24_buffer[clk] = GRF6[24];
    GRF6_25_buffer[clk] = GRF6[25];
    GRF6_26_buffer[clk] = GRF6[26];
    GRF6_27_buffer[clk] = GRF6[27];
    GRF6_28_buffer[clk] = GRF6[28];
    GRF6_29_buffer[clk] = GRF6[29];
    GRF6_30_buffer[clk] = GRF6[30];
    GRF6_31_buffer[clk] = GRF6[31];
    GRF7_0_buffer[clk] = GRF7[0];
    GRF7_1_buffer[clk] = GRF7[1];
    GRF7_2_buffer[clk] = GRF7[2];
    GRF7_3_buffer[clk] = GRF7[3];
    GRF7_4_buffer[clk] = GRF7[4];
    GRF7_5_buffer[clk] = GRF7[5];
    GRF7_6_buffer[clk] = GRF7[6];
    GRF7_7_buffer[clk] = GRF7[7];
    GRF7_8_buffer[clk] = GRF7[8];
    GRF7_9_buffer[clk] = GRF7[9];
    GRF7_10_buffer[clk] = GRF7[10];
    GRF7_11_buffer[clk] = GRF7[11];
    GRF7_12_buffer[clk] = GRF7[12];
    GRF7_13_buffer[clk] = GRF7[13];
    GRF7_14_buffer[clk] = GRF7[14];
    GRF7_15_buffer[clk] = GRF7[15];
    GRF7_16_buffer[clk] = GRF7[16];
    GRF7_17_buffer[clk] = GRF7[17];
    GRF7_18_buffer[clk] = GRF7[18];
    GRF7_19_buffer[clk] = GRF7[19];
    GRF7_20_buffer[clk] = GRF7[20];
    GRF7_21_buffer[clk] = GRF7[21];
    GRF7_22_buffer[clk] = GRF7[22];
    GRF7_23_buffer[clk] = GRF7[23];
    GRF7_24_buffer[clk] = GRF7[24];
    GRF7_25_buffer[clk] = GRF7[25];
    GRF7_26_buffer[clk] = GRF7[26];
    GRF7_27_buffer[clk] = GRF7[27];
    GRF7_28_buffer[clk] = GRF7[28];
    GRF7_29_buffer[clk] = GRF7[29];
    GRF7_30_buffer[clk] = GRF7[30];
    GRF7_31_buffer[clk] = GRF7[31];
    GRF8_0_buffer[clk] = GRF8[0];
    GRF8_1_buffer[clk] = GRF8[1];
    GRF8_2_buffer[clk] = GRF8[2];
    GRF8_3_buffer[clk] = GRF8[3];
    GRF8_4_buffer[clk] = GRF8[4];
    GRF8_5_buffer[clk] = GRF8[5];
    GRF8_6_buffer[clk] = GRF8[6];
    GRF8_7_buffer[clk] = GRF8[7];
    GRF8_8_buffer[clk] = GRF8[8];
    GRF8_9_buffer[clk] = GRF8[9];
    GRF8_10_buffer[clk] = GRF8[10];
    GRF8_11_buffer[clk] = GRF8[11];
    GRF8_12_buffer[clk] = GRF8[12];
    GRF8_13_buffer[clk] = GRF8[13];
    GRF8_14_buffer[clk] = GRF8[14];
    GRF8_15_buffer[clk] = GRF8[15];
    GRF8_16_buffer[clk] = GRF8[16];
    GRF8_17_buffer[clk] = GRF8[17];
    GRF8_18_buffer[clk] = GRF8[18];
    GRF8_19_buffer[clk] = GRF8[19];
    GRF8_20_buffer[clk] = GRF8[20];
    GRF8_21_buffer[clk] = GRF8[21];
    GRF8_22_buffer[clk] = GRF8[22];
    GRF8_23_buffer[clk] = GRF8[23];
    GRF8_24_buffer[clk] = GRF8[24];
    GRF8_25_buffer[clk] = GRF8[25];
    GRF8_26_buffer[clk] = GRF8[26];
    GRF8_27_buffer[clk] = GRF8[27];
    GRF8_28_buffer[clk] = GRF8[28];
    GRF8_29_buffer[clk] = GRF8[29];
    GRF8_30_buffer[clk] = GRF8[30];
    GRF8_31_buffer[clk] = GRF8[31];
    GRF9_0_buffer[clk] = GRF9[0];
    GRF9_1_buffer[clk] = GRF9[1];
    GRF9_2_buffer[clk] = GRF9[2];
    GRF9_3_buffer[clk] = GRF9[3];
    GRF9_4_buffer[clk] = GRF9[4];
    GRF9_5_buffer[clk] = GRF9[5];
    GRF9_6_buffer[clk] = GRF9[6];
    GRF9_7_buffer[clk] = GRF9[7];
    GRF9_8_buffer[clk] = GRF9[8];
    GRF9_9_buffer[clk] = GRF9[9];
    GRF9_10_buffer[clk] = GRF9[10];
    GRF9_11_buffer[clk] = GRF9[11];
    GRF9_12_buffer[clk] = GRF9[12];
    GRF9_13_buffer[clk] = GRF9[13];
    GRF9_14_buffer[clk] = GRF9[14];
    GRF9_15_buffer[clk] = GRF9[15];
    GRF9_16_buffer[clk] = GRF9[16];
    GRF9_17_buffer[clk] = GRF9[17];
    GRF9_18_buffer[clk] = GRF9[18];
    GRF9_19_buffer[clk] = GRF9[19];
    GRF9_20_buffer[clk] = GRF9[20];
    GRF9_21_buffer[clk] = GRF9[21];
    GRF9_22_buffer[clk] = GRF9[22];
    GRF9_23_buffer[clk] = GRF9[23];
    GRF9_24_buffer[clk] = GRF9[24];
    GRF9_25_buffer[clk] = GRF9[25];
    GRF9_26_buffer[clk] = GRF9[26];
    GRF9_27_buffer[clk] = GRF9[27];
    GRF9_28_buffer[clk] = GRF9[28];
    GRF9_29_buffer[clk] = GRF9[29];
    GRF9_30_buffer[clk] = GRF9[30];
    GRF9_31_buffer[clk] = GRF9[31];
    GRF10_0_buffer[clk] = GRF10[0];
    GRF10_1_buffer[clk] = GRF10[1];
    GRF10_2_buffer[clk] = GRF10[2];
    GRF10_3_buffer[clk] = GRF10[3];
    GRF10_4_buffer[clk] = GRF10[4];
    GRF10_5_buffer[clk] = GRF10[5];
    GRF10_6_buffer[clk] = GRF10[6];
    GRF10_7_buffer[clk] = GRF10[7];
    GRF10_8_buffer[clk] = GRF10[8];
    GRF10_9_buffer[clk] = GRF10[9];
    GRF10_10_buffer[clk] = GRF10[10];
    GRF10_11_buffer[clk] = GRF10[11];
    GRF10_12_buffer[clk] = GRF10[12];
    GRF10_13_buffer[clk] = GRF10[13];
    GRF10_14_buffer[clk] = GRF10[14];
    GRF10_15_buffer[clk] = GRF10[15];
    GRF10_16_buffer[clk] = GRF10[16];
    GRF10_17_buffer[clk] = GRF10[17];
    GRF10_18_buffer[clk] = GRF10[18];
    GRF10_19_buffer[clk] = GRF10[19];
    GRF10_20_buffer[clk] = GRF10[20];
    GRF10_21_buffer[clk] = GRF10[21];
    GRF10_22_buffer[clk] = GRF10[22];
    GRF10_23_buffer[clk] = GRF10[23];
    GRF10_24_buffer[clk] = GRF10[24];
    GRF10_25_buffer[clk] = GRF10[25];
    GRF10_26_buffer[clk] = GRF10[26];
    GRF10_27_buffer[clk] = GRF10[27];
    GRF10_28_buffer[clk] = GRF10[28];
    GRF10_29_buffer[clk] = GRF10[29];
    GRF10_30_buffer[clk] = GRF10[30];
    GRF10_31_buffer[clk] = GRF10[31];
    GRF11_0_buffer[clk] = GRF11[0];
    GRF11_1_buffer[clk] = GRF11[1];
    GRF11_2_buffer[clk] = GRF11[2];
    GRF11_3_buffer[clk] = GRF11[3];
    GRF11_4_buffer[clk] = GRF11[4];
    GRF11_5_buffer[clk] = GRF11[5];
    GRF11_6_buffer[clk] = GRF11[6];
    GRF11_7_buffer[clk] = GRF11[7];
    GRF11_8_buffer[clk] = GRF11[8];
    GRF11_9_buffer[clk] = GRF11[9];
    GRF11_10_buffer[clk] = GRF11[10];
    GRF11_11_buffer[clk] = GRF11[11];
    GRF11_12_buffer[clk] = GRF11[12];
    GRF11_13_buffer[clk] = GRF11[13];
    GRF11_14_buffer[clk] = GRF11[14];
    GRF11_15_buffer[clk] = GRF11[15];
    GRF11_16_buffer[clk] = GRF11[16];
    GRF11_17_buffer[clk] = GRF11[17];
    GRF11_18_buffer[clk] = GRF11[18];
    GRF11_19_buffer[clk] = GRF11[19];
    GRF11_20_buffer[clk] = GRF11[20];
    GRF11_21_buffer[clk] = GRF11[21];
    GRF11_22_buffer[clk] = GRF11[22];
    GRF11_23_buffer[clk] = GRF11[23];
    GRF11_24_buffer[clk] = GRF11[24];
    GRF11_25_buffer[clk] = GRF11[25];
    GRF11_26_buffer[clk] = GRF11[26];
    GRF11_27_buffer[clk] = GRF11[27];
    GRF11_28_buffer[clk] = GRF11[28];
    GRF11_29_buffer[clk] = GRF11[29];
    GRF11_30_buffer[clk] = GRF11[30];
    GRF11_31_buffer[clk] = GRF11[31];
    GRF12_0_buffer[clk] = GRF12[0];
    GRF12_1_buffer[clk] = GRF12[1];
    GRF12_2_buffer[clk] = GRF12[2];
    GRF12_3_buffer[clk] = GRF12[3];
    GRF12_4_buffer[clk] = GRF12[4];
    GRF12_5_buffer[clk] = GRF12[5];
    GRF12_6_buffer[clk] = GRF12[6];
    GRF12_7_buffer[clk] = GRF12[7];
    GRF12_8_buffer[clk] = GRF12[8];
    GRF12_9_buffer[clk] = GRF12[9];
    GRF12_10_buffer[clk] = GRF12[10];
    GRF12_11_buffer[clk] = GRF12[11];
    GRF12_12_buffer[clk] = GRF12[12];
    GRF12_13_buffer[clk] = GRF12[13];
    GRF12_14_buffer[clk] = GRF12[14];
    GRF12_15_buffer[clk] = GRF12[15];
    GRF12_16_buffer[clk] = GRF12[16];
    GRF12_17_buffer[clk] = GRF12[17];
    GRF12_18_buffer[clk] = GRF12[18];
    GRF12_19_buffer[clk] = GRF12[19];
    GRF12_20_buffer[clk] = GRF12[20];
    GRF12_21_buffer[clk] = GRF12[21];
    GRF12_22_buffer[clk] = GRF12[22];
    GRF12_23_buffer[clk] = GRF12[23];
    GRF12_24_buffer[clk] = GRF12[24];
    GRF12_25_buffer[clk] = GRF12[25];
    GRF12_26_buffer[clk] = GRF12[26];
    GRF12_27_buffer[clk] = GRF12[27];
    GRF12_28_buffer[clk] = GRF12[28];
    GRF12_29_buffer[clk] = GRF12[29];
    GRF12_30_buffer[clk] = GRF12[30];
    GRF12_31_buffer[clk] = GRF12[31];
    GRF13_0_buffer[clk] = GRF13[0];
    GRF13_1_buffer[clk] = GRF13[1];
    GRF13_2_buffer[clk] = GRF13[2];
    GRF13_3_buffer[clk] = GRF13[3];
    GRF13_4_buffer[clk] = GRF13[4];
    GRF13_5_buffer[clk] = GRF13[5];
    GRF13_6_buffer[clk] = GRF13[6];
    GRF13_7_buffer[clk] = GRF13[7];
    GRF13_8_buffer[clk] = GRF13[8];
    GRF13_9_buffer[clk] = GRF13[9];
    GRF13_10_buffer[clk] = GRF13[10];
    GRF13_11_buffer[clk] = GRF13[11];
    GRF13_12_buffer[clk] = GRF13[12];
    GRF13_13_buffer[clk] = GRF13[13];
    GRF13_14_buffer[clk] = GRF13[14];
    GRF13_15_buffer[clk] = GRF13[15];
    GRF13_16_buffer[clk] = GRF13[16];
    GRF13_17_buffer[clk] = GRF13[17];
    GRF13_18_buffer[clk] = GRF13[18];
    GRF13_19_buffer[clk] = GRF13[19];
    GRF13_20_buffer[clk] = GRF13[20];
    GRF13_21_buffer[clk] = GRF13[21];
    GRF13_22_buffer[clk] = GRF13[22];
    GRF13_23_buffer[clk] = GRF13[23];
    GRF13_24_buffer[clk] = GRF13[24];
    GRF13_25_buffer[clk] = GRF13[25];
    GRF13_26_buffer[clk] = GRF13[26];
    GRF13_27_buffer[clk] = GRF13[27];
    GRF13_28_buffer[clk] = GRF13[28];
    GRF13_29_buffer[clk] = GRF13[29];
    GRF13_30_buffer[clk] = GRF13[30];
    GRF13_31_buffer[clk] = GRF13[31];
    GRF14_0_buffer[clk] = GRF14[0];
    GRF14_1_buffer[clk] = GRF14[1];
    GRF14_2_buffer[clk] = GRF14[2];
    GRF14_3_buffer[clk] = GRF14[3];
    GRF14_4_buffer[clk] = GRF14[4];
    GRF14_5_buffer[clk] = GRF14[5];
    GRF14_6_buffer[clk] = GRF14[6];
    GRF14_7_buffer[clk] = GRF14[7];
    GRF14_8_buffer[clk] = GRF14[8];
    GRF14_9_buffer[clk] = GRF14[9];
    GRF14_10_buffer[clk] = GRF14[10];
    GRF14_11_buffer[clk] = GRF14[11];
    GRF14_12_buffer[clk] = GRF14[12];
    GRF14_13_buffer[clk] = GRF14[13];
    GRF14_14_buffer[clk] = GRF14[14];
    GRF14_15_buffer[clk] = GRF14[15];
    GRF14_16_buffer[clk] = GRF14[16];
    GRF14_17_buffer[clk] = GRF14[17];
    GRF14_18_buffer[clk] = GRF14[18];
    GRF14_19_buffer[clk] = GRF14[19];
    GRF14_20_buffer[clk] = GRF14[20];
    GRF14_21_buffer[clk] = GRF14[21];
    GRF14_22_buffer[clk] = GRF14[22];
    GRF14_23_buffer[clk] = GRF14[23];
    GRF14_24_buffer[clk] = GRF14[24];
    GRF14_25_buffer[clk] = GRF14[25];
    GRF14_26_buffer[clk] = GRF14[26];
    GRF14_27_buffer[clk] = GRF14[27];
    GRF14_28_buffer[clk] = GRF14[28];
    GRF14_29_buffer[clk] = GRF14[29];
    GRF14_30_buffer[clk] = GRF14[30];
    GRF14_31_buffer[clk] = GRF14[31];
    GRF15_0_buffer[clk] = GRF15[0];
    GRF15_1_buffer[clk] = GRF15[1];
    GRF15_2_buffer[clk] = GRF15[2];
    GRF15_3_buffer[clk] = GRF15[3];
    GRF15_4_buffer[clk] = GRF15[4];
    GRF15_5_buffer[clk] = GRF15[5];
    GRF15_6_buffer[clk] = GRF15[6];
    GRF15_7_buffer[clk] = GRF15[7];
    GRF15_8_buffer[clk] = GRF15[8];
    GRF15_9_buffer[clk] = GRF15[9];
    GRF15_10_buffer[clk] = GRF15[10];
    GRF15_11_buffer[clk] = GRF15[11];
    GRF15_12_buffer[clk] = GRF15[12];
    GRF15_13_buffer[clk] = GRF15[13];
    GRF15_14_buffer[clk] = GRF15[14];
    GRF15_15_buffer[clk] = GRF15[15];
    GRF15_16_buffer[clk] = GRF15[16];
    GRF15_17_buffer[clk] = GRF15[17];
    GRF15_18_buffer[clk] = GRF15[18];
    GRF15_19_buffer[clk] = GRF15[19];
    GRF15_20_buffer[clk] = GRF15[20];
    GRF15_21_buffer[clk] = GRF15[21];
    GRF15_22_buffer[clk] = GRF15[22];
    GRF15_23_buffer[clk] = GRF15[23];
    GRF15_24_buffer[clk] = GRF15[24];
    GRF15_25_buffer[clk] = GRF15[25];
    GRF15_26_buffer[clk] = GRF15[26];
    GRF15_27_buffer[clk] = GRF15[27];
    GRF15_28_buffer[clk] = GRF15[28];
    GRF15_29_buffer[clk] = GRF15[29];
    GRF15_30_buffer[clk] = GRF15[30];
    GRF15_31_buffer[clk] = GRF15[31];
    GRF16_0_buffer[clk] = GRF16[0];
    GRF16_1_buffer[clk] = GRF16[1];
    GRF16_2_buffer[clk] = GRF16[2];
    GRF16_3_buffer[clk] = GRF16[3];
    GRF16_4_buffer[clk] = GRF16[4];
    GRF16_5_buffer[clk] = GRF16[5];
    GRF16_6_buffer[clk] = GRF16[6];
    GRF16_7_buffer[clk] = GRF16[7];
    GRF16_8_buffer[clk] = GRF16[8];
    GRF16_9_buffer[clk] = GRF16[9];
    GRF16_10_buffer[clk] = GRF16[10];
    GRF16_11_buffer[clk] = GRF16[11];
    GRF16_12_buffer[clk] = GRF16[12];
    GRF16_13_buffer[clk] = GRF16[13];
    GRF16_14_buffer[clk] = GRF16[14];
    GRF16_15_buffer[clk] = GRF16[15];
    GRF16_16_buffer[clk] = GRF16[16];
    GRF16_17_buffer[clk] = GRF16[17];
    GRF16_18_buffer[clk] = GRF16[18];
    GRF16_19_buffer[clk] = GRF16[19];
    GRF16_20_buffer[clk] = GRF16[20];
    GRF16_21_buffer[clk] = GRF16[21];
    GRF16_22_buffer[clk] = GRF16[22];
    GRF16_23_buffer[clk] = GRF16[23];
    GRF16_24_buffer[clk] = GRF16[24];
    GRF16_25_buffer[clk] = GRF16[25];
    GRF16_26_buffer[clk] = GRF16[26];
    GRF16_27_buffer[clk] = GRF16[27];
    GRF16_28_buffer[clk] = GRF16[28];
    GRF16_29_buffer[clk] = GRF16[29];
    GRF16_30_buffer[clk] = GRF16[30];
    GRF16_31_buffer[clk] = GRF16[31];
    GRF17_0_buffer[clk] = GRF17[0];
    GRF17_1_buffer[clk] = GRF17[1];
    GRF17_2_buffer[clk] = GRF17[2];
    GRF17_3_buffer[clk] = GRF17[3];
    GRF17_4_buffer[clk] = GRF17[4];
    GRF17_5_buffer[clk] = GRF17[5];
    GRF17_6_buffer[clk] = GRF17[6];
    GRF17_7_buffer[clk] = GRF17[7];
    GRF17_8_buffer[clk] = GRF17[8];
    GRF17_9_buffer[clk] = GRF17[9];
    GRF17_10_buffer[clk] = GRF17[10];
    GRF17_11_buffer[clk] = GRF17[11];
    GRF17_12_buffer[clk] = GRF17[12];
    GRF17_13_buffer[clk] = GRF17[13];
    GRF17_14_buffer[clk] = GRF17[14];
    GRF17_15_buffer[clk] = GRF17[15];
    GRF17_16_buffer[clk] = GRF17[16];
    GRF17_17_buffer[clk] = GRF17[17];
    GRF17_18_buffer[clk] = GRF17[18];
    GRF17_19_buffer[clk] = GRF17[19];
    GRF17_20_buffer[clk] = GRF17[20];
    GRF17_21_buffer[clk] = GRF17[21];
    GRF17_22_buffer[clk] = GRF17[22];
    GRF17_23_buffer[clk] = GRF17[23];
    GRF17_24_buffer[clk] = GRF17[24];
    GRF17_25_buffer[clk] = GRF17[25];
    GRF17_26_buffer[clk] = GRF17[26];
    GRF17_27_buffer[clk] = GRF17[27];
    GRF17_28_buffer[clk] = GRF17[28];
    GRF17_29_buffer[clk] = GRF17[29];
    GRF17_30_buffer[clk] = GRF17[30];
    GRF17_31_buffer[clk] = GRF17[31];
    GRF18_0_buffer[clk] = GRF18[0];
    GRF18_1_buffer[clk] = GRF18[1];
    GRF18_2_buffer[clk] = GRF18[2];
    GRF18_3_buffer[clk] = GRF18[3];
    GRF18_4_buffer[clk] = GRF18[4];
    GRF18_5_buffer[clk] = GRF18[5];
    GRF18_6_buffer[clk] = GRF18[6];
    GRF18_7_buffer[clk] = GRF18[7];
    GRF18_8_buffer[clk] = GRF18[8];
    GRF18_9_buffer[clk] = GRF18[9];
    GRF18_10_buffer[clk] = GRF18[10];
    GRF18_11_buffer[clk] = GRF18[11];
    GRF18_12_buffer[clk] = GRF18[12];
    GRF18_13_buffer[clk] = GRF18[13];
    GRF18_14_buffer[clk] = GRF18[14];
    GRF18_15_buffer[clk] = GRF18[15];
    GRF18_16_buffer[clk] = GRF18[16];
    GRF18_17_buffer[clk] = GRF18[17];
    GRF18_18_buffer[clk] = GRF18[18];
    GRF18_19_buffer[clk] = GRF18[19];
    GRF18_20_buffer[clk] = GRF18[20];
    GRF18_21_buffer[clk] = GRF18[21];
    GRF18_22_buffer[clk] = GRF18[22];
    GRF18_23_buffer[clk] = GRF18[23];
    GRF18_24_buffer[clk] = GRF18[24];
    GRF18_25_buffer[clk] = GRF18[25];
    GRF18_26_buffer[clk] = GRF18[26];
    GRF18_27_buffer[clk] = GRF18[27];
    GRF18_28_buffer[clk] = GRF18[28];
    GRF18_29_buffer[clk] = GRF18[29];
    GRF18_30_buffer[clk] = GRF18[30];
    GRF18_31_buffer[clk] = GRF18[31];
    GRF19_0_buffer[clk] = GRF19[0];
    GRF19_1_buffer[clk] = GRF19[1];
    GRF19_2_buffer[clk] = GRF19[2];
    GRF19_3_buffer[clk] = GRF19[3];
    GRF19_4_buffer[clk] = GRF19[4];
    GRF19_5_buffer[clk] = GRF19[5];
    GRF19_6_buffer[clk] = GRF19[6];
    GRF19_7_buffer[clk] = GRF19[7];
    GRF19_8_buffer[clk] = GRF19[8];
    GRF19_9_buffer[clk] = GRF19[9];
    GRF19_10_buffer[clk] = GRF19[10];
    GRF19_11_buffer[clk] = GRF19[11];
    GRF19_12_buffer[clk] = GRF19[12];
    GRF19_13_buffer[clk] = GRF19[13];
    GRF19_14_buffer[clk] = GRF19[14];
    GRF19_15_buffer[clk] = GRF19[15];
    GRF19_16_buffer[clk] = GRF19[16];
    GRF19_17_buffer[clk] = GRF19[17];
    GRF19_18_buffer[clk] = GRF19[18];
    GRF19_19_buffer[clk] = GRF19[19];
    GRF19_20_buffer[clk] = GRF19[20];
    GRF19_21_buffer[clk] = GRF19[21];
    GRF19_22_buffer[clk] = GRF19[22];
    GRF19_23_buffer[clk] = GRF19[23];
    GRF19_24_buffer[clk] = GRF19[24];
    GRF19_25_buffer[clk] = GRF19[25];
    GRF19_26_buffer[clk] = GRF19[26];
    GRF19_27_buffer[clk] = GRF19[27];
    GRF19_28_buffer[clk] = GRF19[28];
    GRF19_29_buffer[clk] = GRF19[29];
    GRF19_30_buffer[clk] = GRF19[30];
    GRF19_31_buffer[clk] = GRF19[31];
    GRF20_0_buffer[clk] = GRF20[0];
    GRF20_1_buffer[clk] = GRF20[1];
    GRF20_2_buffer[clk] = GRF20[2];
    GRF20_3_buffer[clk] = GRF20[3];
    GRF20_4_buffer[clk] = GRF20[4];
    GRF20_5_buffer[clk] = GRF20[5];
    GRF20_6_buffer[clk] = GRF20[6];
    GRF20_7_buffer[clk] = GRF20[7];
    GRF20_8_buffer[clk] = GRF20[8];
    GRF20_9_buffer[clk] = GRF20[9];
    GRF20_10_buffer[clk] = GRF20[10];
    GRF20_11_buffer[clk] = GRF20[11];
    GRF20_12_buffer[clk] = GRF20[12];
    GRF20_13_buffer[clk] = GRF20[13];
    GRF20_14_buffer[clk] = GRF20[14];
    GRF20_15_buffer[clk] = GRF20[15];
    GRF20_16_buffer[clk] = GRF20[16];
    GRF20_17_buffer[clk] = GRF20[17];
    GRF20_18_buffer[clk] = GRF20[18];
    GRF20_19_buffer[clk] = GRF20[19];
    GRF20_20_buffer[clk] = GRF20[20];
    GRF20_21_buffer[clk] = GRF20[21];
    GRF20_22_buffer[clk] = GRF20[22];
    GRF20_23_buffer[clk] = GRF20[23];
    GRF20_24_buffer[clk] = GRF20[24];
    GRF20_25_buffer[clk] = GRF20[25];
    GRF20_26_buffer[clk] = GRF20[26];
    GRF20_27_buffer[clk] = GRF20[27];
    GRF20_28_buffer[clk] = GRF20[28];
    GRF20_29_buffer[clk] = GRF20[29];
    GRF20_30_buffer[clk] = GRF20[30];
    GRF20_31_buffer[clk] = GRF20[31];
    GRF21_0_buffer[clk] = GRF21[0];
    GRF21_1_buffer[clk] = GRF21[1];
    GRF21_2_buffer[clk] = GRF21[2];
    GRF21_3_buffer[clk] = GRF21[3];
    GRF21_4_buffer[clk] = GRF21[4];
    GRF21_5_buffer[clk] = GRF21[5];
    GRF21_6_buffer[clk] = GRF21[6];
    GRF21_7_buffer[clk] = GRF21[7];
    GRF21_8_buffer[clk] = GRF21[8];
    GRF21_9_buffer[clk] = GRF21[9];
    GRF21_10_buffer[clk] = GRF21[10];
    GRF21_11_buffer[clk] = GRF21[11];
    GRF21_12_buffer[clk] = GRF21[12];
    GRF21_13_buffer[clk] = GRF21[13];
    GRF21_14_buffer[clk] = GRF21[14];
    GRF21_15_buffer[clk] = GRF21[15];
    GRF21_16_buffer[clk] = GRF21[16];
    GRF21_17_buffer[clk] = GRF21[17];
    GRF21_18_buffer[clk] = GRF21[18];
    GRF21_19_buffer[clk] = GRF21[19];
    GRF21_20_buffer[clk] = GRF21[20];
    GRF21_21_buffer[clk] = GRF21[21];
    GRF21_22_buffer[clk] = GRF21[22];
    GRF21_23_buffer[clk] = GRF21[23];
    GRF21_24_buffer[clk] = GRF21[24];
    GRF21_25_buffer[clk] = GRF21[25];
    GRF21_26_buffer[clk] = GRF21[26];
    GRF21_27_buffer[clk] = GRF21[27];
    GRF21_28_buffer[clk] = GRF21[28];
    GRF21_29_buffer[clk] = GRF21[29];
    GRF21_30_buffer[clk] = GRF21[30];
    GRF21_31_buffer[clk] = GRF21[31];
    GRF22_0_buffer[clk] = GRF22[0];
    GRF22_1_buffer[clk] = GRF22[1];
    GRF22_2_buffer[clk] = GRF22[2];
    GRF22_3_buffer[clk] = GRF22[3];
    GRF22_4_buffer[clk] = GRF22[4];
    GRF22_5_buffer[clk] = GRF22[5];
    GRF22_6_buffer[clk] = GRF22[6];
    GRF22_7_buffer[clk] = GRF22[7];
    GRF22_8_buffer[clk] = GRF22[8];
    GRF22_9_buffer[clk] = GRF22[9];
    GRF22_10_buffer[clk] = GRF22[10];
    GRF22_11_buffer[clk] = GRF22[11];
    GRF22_12_buffer[clk] = GRF22[12];
    GRF22_13_buffer[clk] = GRF22[13];
    GRF22_14_buffer[clk] = GRF22[14];
    GRF22_15_buffer[clk] = GRF22[15];
    GRF22_16_buffer[clk] = GRF22[16];
    GRF22_17_buffer[clk] = GRF22[17];
    GRF22_18_buffer[clk] = GRF22[18];
    GRF22_19_buffer[clk] = GRF22[19];
    GRF22_20_buffer[clk] = GRF22[20];
    GRF22_21_buffer[clk] = GRF22[21];
    GRF22_22_buffer[clk] = GRF22[22];
    GRF22_23_buffer[clk] = GRF22[23];
    GRF22_24_buffer[clk] = GRF22[24];
    GRF22_25_buffer[clk] = GRF22[25];
    GRF22_26_buffer[clk] = GRF22[26];
    GRF22_27_buffer[clk] = GRF22[27];
    GRF22_28_buffer[clk] = GRF22[28];
    GRF22_29_buffer[clk] = GRF22[29];
    GRF22_30_buffer[clk] = GRF22[30];
    GRF22_31_buffer[clk] = GRF22[31];
    GRF23_0_buffer[clk] = GRF23[0];
    GRF23_1_buffer[clk] = GRF23[1];
    GRF23_2_buffer[clk] = GRF23[2];
    GRF23_3_buffer[clk] = GRF23[3];
    GRF23_4_buffer[clk] = GRF23[4];
    GRF23_5_buffer[clk] = GRF23[5];
    GRF23_6_buffer[clk] = GRF23[6];
    GRF23_7_buffer[clk] = GRF23[7];
    GRF23_8_buffer[clk] = GRF23[8];
    GRF23_9_buffer[clk] = GRF23[9];
    GRF23_10_buffer[clk] = GRF23[10];
    GRF23_11_buffer[clk] = GRF23[11];
    GRF23_12_buffer[clk] = GRF23[12];
    GRF23_13_buffer[clk] = GRF23[13];
    GRF23_14_buffer[clk] = GRF23[14];
    GRF23_15_buffer[clk] = GRF23[15];
    GRF23_16_buffer[clk] = GRF23[16];
    GRF23_17_buffer[clk] = GRF23[17];
    GRF23_18_buffer[clk] = GRF23[18];
    GRF23_19_buffer[clk] = GRF23[19];
    GRF23_20_buffer[clk] = GRF23[20];
    GRF23_21_buffer[clk] = GRF23[21];
    GRF23_22_buffer[clk] = GRF23[22];
    GRF23_23_buffer[clk] = GRF23[23];
    GRF23_24_buffer[clk] = GRF23[24];
    GRF23_25_buffer[clk] = GRF23[25];
    GRF23_26_buffer[clk] = GRF23[26];
    GRF23_27_buffer[clk] = GRF23[27];
    GRF23_28_buffer[clk] = GRF23[28];
    GRF23_29_buffer[clk] = GRF23[29];
    GRF23_30_buffer[clk] = GRF23[30];
    GRF23_31_buffer[clk] = GRF23[31];
    GRF24_0_buffer[clk] = GRF24[0];
    GRF24_1_buffer[clk] = GRF24[1];
    GRF24_2_buffer[clk] = GRF24[2];
    GRF24_3_buffer[clk] = GRF24[3];
    GRF24_4_buffer[clk] = GRF24[4];
    GRF24_5_buffer[clk] = GRF24[5];
    GRF24_6_buffer[clk] = GRF24[6];
    GRF24_7_buffer[clk] = GRF24[7];
    GRF24_8_buffer[clk] = GRF24[8];
    GRF24_9_buffer[clk] = GRF24[9];
    GRF24_10_buffer[clk] = GRF24[10];
    GRF24_11_buffer[clk] = GRF24[11];
    GRF24_12_buffer[clk] = GRF24[12];
    GRF24_13_buffer[clk] = GRF24[13];
    GRF24_14_buffer[clk] = GRF24[14];
    GRF24_15_buffer[clk] = GRF24[15];
    GRF24_16_buffer[clk] = GRF24[16];
    GRF24_17_buffer[clk] = GRF24[17];
    GRF24_18_buffer[clk] = GRF24[18];
    GRF24_19_buffer[clk] = GRF24[19];
    GRF24_20_buffer[clk] = GRF24[20];
    GRF24_21_buffer[clk] = GRF24[21];
    GRF24_22_buffer[clk] = GRF24[22];
    GRF24_23_buffer[clk] = GRF24[23];
    GRF24_24_buffer[clk] = GRF24[24];
    GRF24_25_buffer[clk] = GRF24[25];
    GRF24_26_buffer[clk] = GRF24[26];
    GRF24_27_buffer[clk] = GRF24[27];
    GRF24_28_buffer[clk] = GRF24[28];
    GRF24_29_buffer[clk] = GRF24[29];
    GRF24_30_buffer[clk] = GRF24[30];
    GRF24_31_buffer[clk] = GRF24[31];
    GRF25_0_buffer[clk] = GRF25[0];
    GRF25_1_buffer[clk] = GRF25[1];
    GRF25_2_buffer[clk] = GRF25[2];
    GRF25_3_buffer[clk] = GRF25[3];
    GRF25_4_buffer[clk] = GRF25[4];
    GRF25_5_buffer[clk] = GRF25[5];
    GRF25_6_buffer[clk] = GRF25[6];
    GRF25_7_buffer[clk] = GRF25[7];
    GRF25_8_buffer[clk] = GRF25[8];
    GRF25_9_buffer[clk] = GRF25[9];
    GRF25_10_buffer[clk] = GRF25[10];
    GRF25_11_buffer[clk] = GRF25[11];
    GRF25_12_buffer[clk] = GRF25[12];
    GRF25_13_buffer[clk] = GRF25[13];
    GRF25_14_buffer[clk] = GRF25[14];
    GRF25_15_buffer[clk] = GRF25[15];
    GRF25_16_buffer[clk] = GRF25[16];
    GRF25_17_buffer[clk] = GRF25[17];
    GRF25_18_buffer[clk] = GRF25[18];
    GRF25_19_buffer[clk] = GRF25[19];
    GRF25_20_buffer[clk] = GRF25[20];
    GRF25_21_buffer[clk] = GRF25[21];
    GRF25_22_buffer[clk] = GRF25[22];
    GRF25_23_buffer[clk] = GRF25[23];
    GRF25_24_buffer[clk] = GRF25[24];
    GRF25_25_buffer[clk] = GRF25[25];
    GRF25_26_buffer[clk] = GRF25[26];
    GRF25_27_buffer[clk] = GRF25[27];
    GRF25_28_buffer[clk] = GRF25[28];
    GRF25_29_buffer[clk] = GRF25[29];
    GRF25_30_buffer[clk] = GRF25[30];
    GRF25_31_buffer[clk] = GRF25[31];
    GRF26_0_buffer[clk] = GRF26[0];
    GRF26_1_buffer[clk] = GRF26[1];
    GRF26_2_buffer[clk] = GRF26[2];
    GRF26_3_buffer[clk] = GRF26[3];
    GRF26_4_buffer[clk] = GRF26[4];
    GRF26_5_buffer[clk] = GRF26[5];
    GRF26_6_buffer[clk] = GRF26[6];
    GRF26_7_buffer[clk] = GRF26[7];
    GRF26_8_buffer[clk] = GRF26[8];
    GRF26_9_buffer[clk] = GRF26[9];
    GRF26_10_buffer[clk] = GRF26[10];
    GRF26_11_buffer[clk] = GRF26[11];
    GRF26_12_buffer[clk] = GRF26[12];
    GRF26_13_buffer[clk] = GRF26[13];
    GRF26_14_buffer[clk] = GRF26[14];
    GRF26_15_buffer[clk] = GRF26[15];
    GRF26_16_buffer[clk] = GRF26[16];
    GRF26_17_buffer[clk] = GRF26[17];
    GRF26_18_buffer[clk] = GRF26[18];
    GRF26_19_buffer[clk] = GRF26[19];
    GRF26_20_buffer[clk] = GRF26[20];
    GRF26_21_buffer[clk] = GRF26[21];
    GRF26_22_buffer[clk] = GRF26[22];
    GRF26_23_buffer[clk] = GRF26[23];
    GRF26_24_buffer[clk] = GRF26[24];
    GRF26_25_buffer[clk] = GRF26[25];
    GRF26_26_buffer[clk] = GRF26[26];
    GRF26_27_buffer[clk] = GRF26[27];
    GRF26_28_buffer[clk] = GRF26[28];
    GRF26_29_buffer[clk] = GRF26[29];
    GRF26_30_buffer[clk] = GRF26[30];
    GRF26_31_buffer[clk] = GRF26[31];
    GRF27_0_buffer[clk] = GRF27[0];
    GRF27_1_buffer[clk] = GRF27[1];
    GRF27_2_buffer[clk] = GRF27[2];
    GRF27_3_buffer[clk] = GRF27[3];
    GRF27_4_buffer[clk] = GRF27[4];
    GRF27_5_buffer[clk] = GRF27[5];
    GRF27_6_buffer[clk] = GRF27[6];
    GRF27_7_buffer[clk] = GRF27[7];
    GRF27_8_buffer[clk] = GRF27[8];
    GRF27_9_buffer[clk] = GRF27[9];
    GRF27_10_buffer[clk] = GRF27[10];
    GRF27_11_buffer[clk] = GRF27[11];
    GRF27_12_buffer[clk] = GRF27[12];
    GRF27_13_buffer[clk] = GRF27[13];
    GRF27_14_buffer[clk] = GRF27[14];
    GRF27_15_buffer[clk] = GRF27[15];
    GRF27_16_buffer[clk] = GRF27[16];
    GRF27_17_buffer[clk] = GRF27[17];
    GRF27_18_buffer[clk] = GRF27[18];
    GRF27_19_buffer[clk] = GRF27[19];
    GRF27_20_buffer[clk] = GRF27[20];
    GRF27_21_buffer[clk] = GRF27[21];
    GRF27_22_buffer[clk] = GRF27[22];
    GRF27_23_buffer[clk] = GRF27[23];
    GRF27_24_buffer[clk] = GRF27[24];
    GRF27_25_buffer[clk] = GRF27[25];
    GRF27_26_buffer[clk] = GRF27[26];
    GRF27_27_buffer[clk] = GRF27[27];
    GRF27_28_buffer[clk] = GRF27[28];
    GRF27_29_buffer[clk] = GRF27[29];
    GRF27_30_buffer[clk] = GRF27[30];
    GRF27_31_buffer[clk] = GRF27[31];
    GRF28_0_buffer[clk] = GRF28[0];
    GRF28_1_buffer[clk] = GRF28[1];
    GRF28_2_buffer[clk] = GRF28[2];
    GRF28_3_buffer[clk] = GRF28[3];
    GRF28_4_buffer[clk] = GRF28[4];
    GRF28_5_buffer[clk] = GRF28[5];
    GRF28_6_buffer[clk] = GRF28[6];
    GRF28_7_buffer[clk] = GRF28[7];
    GRF28_8_buffer[clk] = GRF28[8];
    GRF28_9_buffer[clk] = GRF28[9];
    GRF28_10_buffer[clk] = GRF28[10];
    GRF28_11_buffer[clk] = GRF28[11];
    GRF28_12_buffer[clk] = GRF28[12];
    GRF28_13_buffer[clk] = GRF28[13];
    GRF28_14_buffer[clk] = GRF28[14];
    GRF28_15_buffer[clk] = GRF28[15];
    GRF28_16_buffer[clk] = GRF28[16];
    GRF28_17_buffer[clk] = GRF28[17];
    GRF28_18_buffer[clk] = GRF28[18];
    GRF28_19_buffer[clk] = GRF28[19];
    GRF28_20_buffer[clk] = GRF28[20];
    GRF28_21_buffer[clk] = GRF28[21];
    GRF28_22_buffer[clk] = GRF28[22];
    GRF28_23_buffer[clk] = GRF28[23];
    GRF28_24_buffer[clk] = GRF28[24];
    GRF28_25_buffer[clk] = GRF28[25];
    GRF28_26_buffer[clk] = GRF28[26];
    GRF28_27_buffer[clk] = GRF28[27];
    GRF28_28_buffer[clk] = GRF28[28];
    GRF28_29_buffer[clk] = GRF28[29];
    GRF28_30_buffer[clk] = GRF28[30];
    GRF28_31_buffer[clk] = GRF28[31];
    GRF29_0_buffer[clk] = GRF29[0];
    GRF29_1_buffer[clk] = GRF29[1];
    GRF29_2_buffer[clk] = GRF29[2];
    GRF29_3_buffer[clk] = GRF29[3];
    GRF29_4_buffer[clk] = GRF29[4];
    GRF29_5_buffer[clk] = GRF29[5];
    GRF29_6_buffer[clk] = GRF29[6];
    GRF29_7_buffer[clk] = GRF29[7];
    GRF29_8_buffer[clk] = GRF29[8];
    GRF29_9_buffer[clk] = GRF29[9];
    GRF29_10_buffer[clk] = GRF29[10];
    GRF29_11_buffer[clk] = GRF29[11];
    GRF29_12_buffer[clk] = GRF29[12];
    GRF29_13_buffer[clk] = GRF29[13];
    GRF29_14_buffer[clk] = GRF29[14];
    GRF29_15_buffer[clk] = GRF29[15];
    GRF29_16_buffer[clk] = GRF29[16];
    GRF29_17_buffer[clk] = GRF29[17];
    GRF29_18_buffer[clk] = GRF29[18];
    GRF29_19_buffer[clk] = GRF29[19];
    GRF29_20_buffer[clk] = GRF29[20];
    GRF29_21_buffer[clk] = GRF29[21];
    GRF29_22_buffer[clk] = GRF29[22];
    GRF29_23_buffer[clk] = GRF29[23];
    GRF29_24_buffer[clk] = GRF29[24];
    GRF29_25_buffer[clk] = GRF29[25];
    GRF29_26_buffer[clk] = GRF29[26];
    GRF29_27_buffer[clk] = GRF29[27];
    GRF29_28_buffer[clk] = GRF29[28];
    GRF29_29_buffer[clk] = GRF29[29];
    GRF29_30_buffer[clk] = GRF29[30];
    GRF29_31_buffer[clk] = GRF29[31];
    GRF30_0_buffer[clk] = GRF30[0];
    GRF30_1_buffer[clk] = GRF30[1];
    GRF30_2_buffer[clk] = GRF30[2];
    GRF30_3_buffer[clk] = GRF30[3];
    GRF30_4_buffer[clk] = GRF30[4];
    GRF30_5_buffer[clk] = GRF30[5];
    GRF30_6_buffer[clk] = GRF30[6];
    GRF30_7_buffer[clk] = GRF30[7];
    GRF30_8_buffer[clk] = GRF30[8];
    GRF30_9_buffer[clk] = GRF30[9];
    GRF30_10_buffer[clk] = GRF30[10];
    GRF30_11_buffer[clk] = GRF30[11];
    GRF30_12_buffer[clk] = GRF30[12];
    GRF30_13_buffer[clk] = GRF30[13];
    GRF30_14_buffer[clk] = GRF30[14];
    GRF30_15_buffer[clk] = GRF30[15];
    GRF30_16_buffer[clk] = GRF30[16];
    GRF30_17_buffer[clk] = GRF30[17];
    GRF30_18_buffer[clk] = GRF30[18];
    GRF30_19_buffer[clk] = GRF30[19];
    GRF30_20_buffer[clk] = GRF30[20];
    GRF30_21_buffer[clk] = GRF30[21];
    GRF30_22_buffer[clk] = GRF30[22];
    GRF30_23_buffer[clk] = GRF30[23];
    GRF30_24_buffer[clk] = GRF30[24];
    GRF30_25_buffer[clk] = GRF30[25];
    GRF30_26_buffer[clk] = GRF30[26];
    GRF30_27_buffer[clk] = GRF30[27];
    GRF30_28_buffer[clk] = GRF30[28];
    GRF30_29_buffer[clk] = GRF30[29];
    GRF30_30_buffer[clk] = GRF30[30];
    GRF30_31_buffer[clk] = GRF30[31];
    GRF31_0_buffer[clk] = GRF31[0];
    GRF31_1_buffer[clk] = GRF31[1];
    GRF31_2_buffer[clk] = GRF31[2];
    GRF31_3_buffer[clk] = GRF31[3];
    GRF31_4_buffer[clk] = GRF31[4];
    GRF31_5_buffer[clk] = GRF31[5];
    GRF31_6_buffer[clk] = GRF31[6];
    GRF31_7_buffer[clk] = GRF31[7];
    GRF31_8_buffer[clk] = GRF31[8];
    GRF31_9_buffer[clk] = GRF31[9];
    GRF31_10_buffer[clk] = GRF31[10];
    GRF31_11_buffer[clk] = GRF31[11];
    GRF31_12_buffer[clk] = GRF31[12];
    GRF31_13_buffer[clk] = GRF31[13];
    GRF31_14_buffer[clk] = GRF31[14];
    GRF31_15_buffer[clk] = GRF31[15];
    GRF31_16_buffer[clk] = GRF31[16];
    GRF31_17_buffer[clk] = GRF31[17];
    GRF31_18_buffer[clk] = GRF31[18];
    GRF31_19_buffer[clk] = GRF31[19];
    GRF31_20_buffer[clk] = GRF31[20];
    GRF31_21_buffer[clk] = GRF31[21];
    GRF31_22_buffer[clk] = GRF31[22];
    GRF31_23_buffer[clk] = GRF31[23];
    GRF31_24_buffer[clk] = GRF31[24];
    GRF31_25_buffer[clk] = GRF31[25];
    GRF31_26_buffer[clk] = GRF31[26];
    GRF31_27_buffer[clk] = GRF31[27];
    GRF31_28_buffer[clk] = GRF31[28];
    GRF31_29_buffer[clk] = GRF31[29];
    GRF31_30_buffer[clk] = GRF31[30];
    GRF31_31_buffer[clk] = GRF31[31];
    GRF32_0_buffer[clk] = GRF32[0];
    GRF32_1_buffer[clk] = GRF32[1];
    GRF32_2_buffer[clk] = GRF32[2];
    GRF32_3_buffer[clk] = GRF32[3];
    GRF32_4_buffer[clk] = GRF32[4];
    GRF32_5_buffer[clk] = GRF32[5];
    GRF32_6_buffer[clk] = GRF32[6];
    GRF32_7_buffer[clk] = GRF32[7];
    GRF32_8_buffer[clk] = GRF32[8];
    GRF32_9_buffer[clk] = GRF32[9];
    GRF32_10_buffer[clk] = GRF32[10];
    GRF32_11_buffer[clk] = GRF32[11];
    GRF32_12_buffer[clk] = GRF32[12];
    GRF32_13_buffer[clk] = GRF32[13];
    GRF32_14_buffer[clk] = GRF32[14];
    GRF32_15_buffer[clk] = GRF32[15];
    GRF32_16_buffer[clk] = GRF32[16];
    GRF32_17_buffer[clk] = GRF32[17];
    GRF32_18_buffer[clk] = GRF32[18];
    GRF32_19_buffer[clk] = GRF32[19];
    GRF32_20_buffer[clk] = GRF32[20];
    GRF32_21_buffer[clk] = GRF32[21];
    GRF32_22_buffer[clk] = GRF32[22];
    GRF32_23_buffer[clk] = GRF32[23];
    GRF32_24_buffer[clk] = GRF32[24];
    GRF32_25_buffer[clk] = GRF32[25];
    GRF32_26_buffer[clk] = GRF32[26];
    GRF32_27_buffer[clk] = GRF32[27];
    GRF32_28_buffer[clk] = GRF32[28];
    GRF32_29_buffer[clk] = GRF32[29];
    GRF32_30_buffer[clk] = GRF32[30];
    GRF32_31_buffer[clk] = GRF32[31];
    GRF33_0_buffer[clk] = GRF33[0];
    GRF33_1_buffer[clk] = GRF33[1];
    GRF33_2_buffer[clk] = GRF33[2];
    GRF33_3_buffer[clk] = GRF33[3];
    GRF33_4_buffer[clk] = GRF33[4];
    GRF33_5_buffer[clk] = GRF33[5];
    GRF33_6_buffer[clk] = GRF33[6];
    GRF33_7_buffer[clk] = GRF33[7];
    GRF33_8_buffer[clk] = GRF33[8];
    GRF33_9_buffer[clk] = GRF33[9];
    GRF33_10_buffer[clk] = GRF33[10];
    GRF33_11_buffer[clk] = GRF33[11];
    GRF33_12_buffer[clk] = GRF33[12];
    GRF33_13_buffer[clk] = GRF33[13];
    GRF33_14_buffer[clk] = GRF33[14];
    GRF33_15_buffer[clk] = GRF33[15];
    GRF33_16_buffer[clk] = GRF33[16];
    GRF33_17_buffer[clk] = GRF33[17];
    GRF33_18_buffer[clk] = GRF33[18];
    GRF33_19_buffer[clk] = GRF33[19];
    GRF33_20_buffer[clk] = GRF33[20];
    GRF33_21_buffer[clk] = GRF33[21];
    GRF33_22_buffer[clk] = GRF33[22];
    GRF33_23_buffer[clk] = GRF33[23];
    GRF33_24_buffer[clk] = GRF33[24];
    GRF33_25_buffer[clk] = GRF33[25];
    GRF33_26_buffer[clk] = GRF33[26];
    GRF33_27_buffer[clk] = GRF33[27];
    GRF33_28_buffer[clk] = GRF33[28];
    GRF33_29_buffer[clk] = GRF33[29];
    GRF33_30_buffer[clk] = GRF33[30];
    GRF33_31_buffer[clk] = GRF33[31];
    GRF34_0_buffer[clk] = GRF34[0];
    GRF34_1_buffer[clk] = GRF34[1];
    GRF34_2_buffer[clk] = GRF34[2];
    GRF34_3_buffer[clk] = GRF34[3];
    GRF34_4_buffer[clk] = GRF34[4];
    GRF34_5_buffer[clk] = GRF34[5];
    GRF34_6_buffer[clk] = GRF34[6];
    GRF34_7_buffer[clk] = GRF34[7];
    GRF34_8_buffer[clk] = GRF34[8];
    GRF34_9_buffer[clk] = GRF34[9];
    GRF34_10_buffer[clk] = GRF34[10];
    GRF34_11_buffer[clk] = GRF34[11];
    GRF34_12_buffer[clk] = GRF34[12];
    GRF34_13_buffer[clk] = GRF34[13];
    GRF34_14_buffer[clk] = GRF34[14];
    GRF34_15_buffer[clk] = GRF34[15];
    GRF34_16_buffer[clk] = GRF34[16];
    GRF34_17_buffer[clk] = GRF34[17];
    GRF34_18_buffer[clk] = GRF34[18];
    GRF34_19_buffer[clk] = GRF34[19];
    GRF34_20_buffer[clk] = GRF34[20];
    GRF34_21_buffer[clk] = GRF34[21];
    GRF34_22_buffer[clk] = GRF34[22];
    GRF34_23_buffer[clk] = GRF34[23];
    GRF34_24_buffer[clk] = GRF34[24];
    GRF34_25_buffer[clk] = GRF34[25];
    GRF34_26_buffer[clk] = GRF34[26];
    GRF34_27_buffer[clk] = GRF34[27];
    GRF34_28_buffer[clk] = GRF34[28];
    GRF34_29_buffer[clk] = GRF34[29];
    GRF34_30_buffer[clk] = GRF34[30];
    GRF34_31_buffer[clk] = GRF34[31];
    GRF35_0_buffer[clk] = GRF35[0];
    GRF35_1_buffer[clk] = GRF35[1];
    GRF35_2_buffer[clk] = GRF35[2];
    GRF35_3_buffer[clk] = GRF35[3];
    GRF35_4_buffer[clk] = GRF35[4];
    GRF35_5_buffer[clk] = GRF35[5];
    GRF35_6_buffer[clk] = GRF35[6];
    GRF35_7_buffer[clk] = GRF35[7];
    GRF35_8_buffer[clk] = GRF35[8];
    GRF35_9_buffer[clk] = GRF35[9];
    GRF35_10_buffer[clk] = GRF35[10];
    GRF35_11_buffer[clk] = GRF35[11];
    GRF35_12_buffer[clk] = GRF35[12];
    GRF35_13_buffer[clk] = GRF35[13];
    GRF35_14_buffer[clk] = GRF35[14];
    GRF35_15_buffer[clk] = GRF35[15];
    GRF35_16_buffer[clk] = GRF35[16];
    GRF35_17_buffer[clk] = GRF35[17];
    GRF35_18_buffer[clk] = GRF35[18];
    GRF35_19_buffer[clk] = GRF35[19];
    GRF35_20_buffer[clk] = GRF35[20];
    GRF35_21_buffer[clk] = GRF35[21];
    GRF35_22_buffer[clk] = GRF35[22];
    GRF35_23_buffer[clk] = GRF35[23];
    GRF35_24_buffer[clk] = GRF35[24];
    GRF35_25_buffer[clk] = GRF35[25];
    GRF35_26_buffer[clk] = GRF35[26];
    GRF35_27_buffer[clk] = GRF35[27];
    GRF35_28_buffer[clk] = GRF35[28];
    GRF35_29_buffer[clk] = GRF35[29];
    GRF35_30_buffer[clk] = GRF35[30];
    GRF35_31_buffer[clk] = GRF35[31];
    GRF36_0_buffer[clk] = GRF36[0];
    GRF36_1_buffer[clk] = GRF36[1];
    GRF36_2_buffer[clk] = GRF36[2];
    GRF36_3_buffer[clk] = GRF36[3];
    GRF36_4_buffer[clk] = GRF36[4];
    GRF36_5_buffer[clk] = GRF36[5];
    GRF36_6_buffer[clk] = GRF36[6];
    GRF36_7_buffer[clk] = GRF36[7];
    GRF36_8_buffer[clk] = GRF36[8];
    GRF36_9_buffer[clk] = GRF36[9];
    GRF36_10_buffer[clk] = GRF36[10];
    GRF36_11_buffer[clk] = GRF36[11];
    GRF36_12_buffer[clk] = GRF36[12];
    GRF36_13_buffer[clk] = GRF36[13];
    GRF36_14_buffer[clk] = GRF36[14];
    GRF36_15_buffer[clk] = GRF36[15];
    GRF36_16_buffer[clk] = GRF36[16];
    GRF36_17_buffer[clk] = GRF36[17];
    GRF36_18_buffer[clk] = GRF36[18];
    GRF36_19_buffer[clk] = GRF36[19];
    GRF36_20_buffer[clk] = GRF36[20];
    GRF36_21_buffer[clk] = GRF36[21];
    GRF36_22_buffer[clk] = GRF36[22];
    GRF36_23_buffer[clk] = GRF36[23];
    GRF36_24_buffer[clk] = GRF36[24];
    GRF36_25_buffer[clk] = GRF36[25];
    GRF36_26_buffer[clk] = GRF36[26];
    GRF36_27_buffer[clk] = GRF36[27];
    GRF36_28_buffer[clk] = GRF36[28];
    GRF36_29_buffer[clk] = GRF36[29];
    GRF36_30_buffer[clk] = GRF36[30];
    GRF36_31_buffer[clk] = GRF36[31];
    GRF37_0_buffer[clk] = GRF37[0];
    GRF37_1_buffer[clk] = GRF37[1];
    GRF37_2_buffer[clk] = GRF37[2];
    GRF37_3_buffer[clk] = GRF37[3];
    GRF37_4_buffer[clk] = GRF37[4];
    GRF37_5_buffer[clk] = GRF37[5];
    GRF37_6_buffer[clk] = GRF37[6];
    GRF37_7_buffer[clk] = GRF37[7];
    GRF37_8_buffer[clk] = GRF37[8];
    GRF37_9_buffer[clk] = GRF37[9];
    GRF37_10_buffer[clk] = GRF37[10];
    GRF37_11_buffer[clk] = GRF37[11];
    GRF37_12_buffer[clk] = GRF37[12];
    GRF37_13_buffer[clk] = GRF37[13];
    GRF37_14_buffer[clk] = GRF37[14];
    GRF37_15_buffer[clk] = GRF37[15];
    GRF37_16_buffer[clk] = GRF37[16];
    GRF37_17_buffer[clk] = GRF37[17];
    GRF37_18_buffer[clk] = GRF37[18];
    GRF37_19_buffer[clk] = GRF37[19];
    GRF37_20_buffer[clk] = GRF37[20];
    GRF37_21_buffer[clk] = GRF37[21];
    GRF37_22_buffer[clk] = GRF37[22];
    GRF37_23_buffer[clk] = GRF37[23];
    GRF37_24_buffer[clk] = GRF37[24];
    GRF37_25_buffer[clk] = GRF37[25];
    GRF37_26_buffer[clk] = GRF37[26];
    GRF37_27_buffer[clk] = GRF37[27];
    GRF37_28_buffer[clk] = GRF37[28];
    GRF37_29_buffer[clk] = GRF37[29];
    GRF37_30_buffer[clk] = GRF37[30];
    GRF37_31_buffer[clk] = GRF37[31];
    GRF38_0_buffer[clk] = GRF38[0];
    GRF38_1_buffer[clk] = GRF38[1];
    GRF38_2_buffer[clk] = GRF38[2];
    GRF38_3_buffer[clk] = GRF38[3];
    GRF38_4_buffer[clk] = GRF38[4];
    GRF38_5_buffer[clk] = GRF38[5];
    GRF38_6_buffer[clk] = GRF38[6];
    GRF38_7_buffer[clk] = GRF38[7];
    GRF38_8_buffer[clk] = GRF38[8];
    GRF38_9_buffer[clk] = GRF38[9];
    GRF38_10_buffer[clk] = GRF38[10];
    GRF38_11_buffer[clk] = GRF38[11];
    GRF38_12_buffer[clk] = GRF38[12];
    GRF38_13_buffer[clk] = GRF38[13];
    GRF38_14_buffer[clk] = GRF38[14];
    GRF38_15_buffer[clk] = GRF38[15];
    GRF38_16_buffer[clk] = GRF38[16];
    GRF38_17_buffer[clk] = GRF38[17];
    GRF38_18_buffer[clk] = GRF38[18];
    GRF38_19_buffer[clk] = GRF38[19];
    GRF38_20_buffer[clk] = GRF38[20];
    GRF38_21_buffer[clk] = GRF38[21];
    GRF38_22_buffer[clk] = GRF38[22];
    GRF38_23_buffer[clk] = GRF38[23];
    GRF38_24_buffer[clk] = GRF38[24];
    GRF38_25_buffer[clk] = GRF38[25];
    GRF38_26_buffer[clk] = GRF38[26];
    GRF38_27_buffer[clk] = GRF38[27];
    GRF38_28_buffer[clk] = GRF38[28];
    GRF38_29_buffer[clk] = GRF38[29];
    GRF38_30_buffer[clk] = GRF38[30];
    GRF38_31_buffer[clk] = GRF38[31];
    GRF39_0_buffer[clk] = GRF39[0];
    GRF39_1_buffer[clk] = GRF39[1];
    GRF39_2_buffer[clk] = GRF39[2];
    GRF39_3_buffer[clk] = GRF39[3];
    GRF39_4_buffer[clk] = GRF39[4];
    GRF39_5_buffer[clk] = GRF39[5];
    GRF39_6_buffer[clk] = GRF39[6];
    GRF39_7_buffer[clk] = GRF39[7];
    GRF39_8_buffer[clk] = GRF39[8];
    GRF39_9_buffer[clk] = GRF39[9];
    GRF39_10_buffer[clk] = GRF39[10];
    GRF39_11_buffer[clk] = GRF39[11];
    GRF39_12_buffer[clk] = GRF39[12];
    GRF39_13_buffer[clk] = GRF39[13];
    GRF39_14_buffer[clk] = GRF39[14];
    GRF39_15_buffer[clk] = GRF39[15];
    GRF39_16_buffer[clk] = GRF39[16];
    GRF39_17_buffer[clk] = GRF39[17];
    GRF39_18_buffer[clk] = GRF39[18];
    GRF39_19_buffer[clk] = GRF39[19];
    GRF39_20_buffer[clk] = GRF39[20];
    GRF39_21_buffer[clk] = GRF39[21];
    GRF39_22_buffer[clk] = GRF39[22];
    GRF39_23_buffer[clk] = GRF39[23];
    GRF39_24_buffer[clk] = GRF39[24];
    GRF39_25_buffer[clk] = GRF39[25];
    GRF39_26_buffer[clk] = GRF39[26];
    GRF39_27_buffer[clk] = GRF39[27];
    GRF39_28_buffer[clk] = GRF39[28];
    GRF39_29_buffer[clk] = GRF39[29];
    GRF39_30_buffer[clk] = GRF39[30];
    GRF39_31_buffer[clk] = GRF39[31];
    GRF40_0_buffer[clk] = GRF40[0];
    GRF40_1_buffer[clk] = GRF40[1];
    GRF40_2_buffer[clk] = GRF40[2];
    GRF40_3_buffer[clk] = GRF40[3];
    GRF40_4_buffer[clk] = GRF40[4];
    GRF40_5_buffer[clk] = GRF40[5];
    GRF40_6_buffer[clk] = GRF40[6];
    GRF40_7_buffer[clk] = GRF40[7];
    GRF40_8_buffer[clk] = GRF40[8];
    GRF40_9_buffer[clk] = GRF40[9];
    GRF40_10_buffer[clk] = GRF40[10];
    GRF40_11_buffer[clk] = GRF40[11];
    GRF40_12_buffer[clk] = GRF40[12];
    GRF40_13_buffer[clk] = GRF40[13];
    GRF40_14_buffer[clk] = GRF40[14];
    GRF40_15_buffer[clk] = GRF40[15];
    GRF40_16_buffer[clk] = GRF40[16];
    GRF40_17_buffer[clk] = GRF40[17];
    GRF40_18_buffer[clk] = GRF40[18];
    GRF40_19_buffer[clk] = GRF40[19];
    GRF40_20_buffer[clk] = GRF40[20];
    GRF40_21_buffer[clk] = GRF40[21];
    GRF40_22_buffer[clk] = GRF40[22];
    GRF40_23_buffer[clk] = GRF40[23];
    GRF40_24_buffer[clk] = GRF40[24];
    GRF40_25_buffer[clk] = GRF40[25];
    GRF40_26_buffer[clk] = GRF40[26];
    GRF40_27_buffer[clk] = GRF40[27];
    GRF40_28_buffer[clk] = GRF40[28];
    GRF40_29_buffer[clk] = GRF40[29];
    GRF40_30_buffer[clk] = GRF40[30];
    GRF40_31_buffer[clk] = GRF40[31];
    GRF41_0_buffer[clk] = GRF41[0];
    GRF41_1_buffer[clk] = GRF41[1];
    GRF41_2_buffer[clk] = GRF41[2];
    GRF41_3_buffer[clk] = GRF41[3];
    GRF41_4_buffer[clk] = GRF41[4];
    GRF41_5_buffer[clk] = GRF41[5];
    GRF41_6_buffer[clk] = GRF41[6];
    GRF41_7_buffer[clk] = GRF41[7];
    GRF41_8_buffer[clk] = GRF41[8];
    GRF41_9_buffer[clk] = GRF41[9];
    GRF41_10_buffer[clk] = GRF41[10];
    GRF41_11_buffer[clk] = GRF41[11];
    GRF41_12_buffer[clk] = GRF41[12];
    GRF41_13_buffer[clk] = GRF41[13];
    GRF41_14_buffer[clk] = GRF41[14];
    GRF41_15_buffer[clk] = GRF41[15];
    GRF41_16_buffer[clk] = GRF41[16];
    GRF41_17_buffer[clk] = GRF41[17];
    GRF41_18_buffer[clk] = GRF41[18];
    GRF41_19_buffer[clk] = GRF41[19];
    GRF41_20_buffer[clk] = GRF41[20];
    GRF41_21_buffer[clk] = GRF41[21];
    GRF41_22_buffer[clk] = GRF41[22];
    GRF41_23_buffer[clk] = GRF41[23];
    GRF41_24_buffer[clk] = GRF41[24];
    GRF41_25_buffer[clk] = GRF41[25];
    GRF41_26_buffer[clk] = GRF41[26];
    GRF41_27_buffer[clk] = GRF41[27];
    GRF41_28_buffer[clk] = GRF41[28];
    GRF41_29_buffer[clk] = GRF41[29];
    GRF41_30_buffer[clk] = GRF41[30];
    GRF41_31_buffer[clk] = GRF41[31];
    GRF42_0_buffer[clk] = GRF42[0];
    GRF42_1_buffer[clk] = GRF42[1];
    GRF42_2_buffer[clk] = GRF42[2];
    GRF42_3_buffer[clk] = GRF42[3];
    GRF42_4_buffer[clk] = GRF42[4];
    GRF42_5_buffer[clk] = GRF42[5];
    GRF42_6_buffer[clk] = GRF42[6];
    GRF42_7_buffer[clk] = GRF42[7];
    GRF42_8_buffer[clk] = GRF42[8];
    GRF42_9_buffer[clk] = GRF42[9];
    GRF42_10_buffer[clk] = GRF42[10];
    GRF42_11_buffer[clk] = GRF42[11];
    GRF42_12_buffer[clk] = GRF42[12];
    GRF42_13_buffer[clk] = GRF42[13];
    GRF42_14_buffer[clk] = GRF42[14];
    GRF42_15_buffer[clk] = GRF42[15];
    GRF42_16_buffer[clk] = GRF42[16];
    GRF42_17_buffer[clk] = GRF42[17];
    GRF42_18_buffer[clk] = GRF42[18];
    GRF42_19_buffer[clk] = GRF42[19];
    GRF42_20_buffer[clk] = GRF42[20];
    GRF42_21_buffer[clk] = GRF42[21];
    GRF42_22_buffer[clk] = GRF42[22];
    GRF42_23_buffer[clk] = GRF42[23];
    GRF42_24_buffer[clk] = GRF42[24];
    GRF42_25_buffer[clk] = GRF42[25];
    GRF42_26_buffer[clk] = GRF42[26];
    GRF42_27_buffer[clk] = GRF42[27];
    GRF42_28_buffer[clk] = GRF42[28];
    GRF42_29_buffer[clk] = GRF42[29];
    GRF42_30_buffer[clk] = GRF42[30];
    GRF42_31_buffer[clk] = GRF42[31];
    GRF43_0_buffer[clk] = GRF43[0];
    GRF43_1_buffer[clk] = GRF43[1];
    GRF43_2_buffer[clk] = GRF43[2];
    GRF43_3_buffer[clk] = GRF43[3];
    GRF43_4_buffer[clk] = GRF43[4];
    GRF43_5_buffer[clk] = GRF43[5];
    GRF43_6_buffer[clk] = GRF43[6];
    GRF43_7_buffer[clk] = GRF43[7];
    GRF43_8_buffer[clk] = GRF43[8];
    GRF43_9_buffer[clk] = GRF43[9];
    GRF43_10_buffer[clk] = GRF43[10];
    GRF43_11_buffer[clk] = GRF43[11];
    GRF43_12_buffer[clk] = GRF43[12];
    GRF43_13_buffer[clk] = GRF43[13];
    GRF43_14_buffer[clk] = GRF43[14];
    GRF43_15_buffer[clk] = GRF43[15];
    GRF43_16_buffer[clk] = GRF43[16];
    GRF43_17_buffer[clk] = GRF43[17];
    GRF43_18_buffer[clk] = GRF43[18];
    GRF43_19_buffer[clk] = GRF43[19];
    GRF43_20_buffer[clk] = GRF43[20];
    GRF43_21_buffer[clk] = GRF43[21];
    GRF43_22_buffer[clk] = GRF43[22];
    GRF43_23_buffer[clk] = GRF43[23];
    GRF43_24_buffer[clk] = GRF43[24];
    GRF43_25_buffer[clk] = GRF43[25];
    GRF43_26_buffer[clk] = GRF43[26];
    GRF43_27_buffer[clk] = GRF43[27];
    GRF43_28_buffer[clk] = GRF43[28];
    GRF43_29_buffer[clk] = GRF43[29];
    GRF43_30_buffer[clk] = GRF43[30];
    GRF43_31_buffer[clk] = GRF43[31];
    GRF44_0_buffer[clk] = GRF44[0];
    GRF44_1_buffer[clk] = GRF44[1];
    GRF44_2_buffer[clk] = GRF44[2];
    GRF44_3_buffer[clk] = GRF44[3];
    GRF44_4_buffer[clk] = GRF44[4];
    GRF44_5_buffer[clk] = GRF44[5];
    GRF44_6_buffer[clk] = GRF44[6];
    GRF44_7_buffer[clk] = GRF44[7];
    GRF44_8_buffer[clk] = GRF44[8];
    GRF44_9_buffer[clk] = GRF44[9];
    GRF44_10_buffer[clk] = GRF44[10];
    GRF44_11_buffer[clk] = GRF44[11];
    GRF44_12_buffer[clk] = GRF44[12];
    GRF44_13_buffer[clk] = GRF44[13];
    GRF44_14_buffer[clk] = GRF44[14];
    GRF44_15_buffer[clk] = GRF44[15];
    GRF44_16_buffer[clk] = GRF44[16];
    GRF44_17_buffer[clk] = GRF44[17];
    GRF44_18_buffer[clk] = GRF44[18];
    GRF44_19_buffer[clk] = GRF44[19];
    GRF44_20_buffer[clk] = GRF44[20];
    GRF44_21_buffer[clk] = GRF44[21];
    GRF44_22_buffer[clk] = GRF44[22];
    GRF44_23_buffer[clk] = GRF44[23];
    GRF44_24_buffer[clk] = GRF44[24];
    GRF44_25_buffer[clk] = GRF44[25];
    GRF44_26_buffer[clk] = GRF44[26];
    GRF44_27_buffer[clk] = GRF44[27];
    GRF44_28_buffer[clk] = GRF44[28];
    GRF44_29_buffer[clk] = GRF44[29];
    GRF44_30_buffer[clk] = GRF44[30];
    GRF44_31_buffer[clk] = GRF44[31];
    GRF45_0_buffer[clk] = GRF45[0];
    GRF45_1_buffer[clk] = GRF45[1];
    GRF45_2_buffer[clk] = GRF45[2];
    GRF45_3_buffer[clk] = GRF45[3];
    GRF45_4_buffer[clk] = GRF45[4];
    GRF45_5_buffer[clk] = GRF45[5];
    GRF45_6_buffer[clk] = GRF45[6];
    GRF45_7_buffer[clk] = GRF45[7];
    GRF45_8_buffer[clk] = GRF45[8];
    GRF45_9_buffer[clk] = GRF45[9];
    GRF45_10_buffer[clk] = GRF45[10];
    GRF45_11_buffer[clk] = GRF45[11];
    GRF45_12_buffer[clk] = GRF45[12];
    GRF45_13_buffer[clk] = GRF45[13];
    GRF45_14_buffer[clk] = GRF45[14];
    GRF45_15_buffer[clk] = GRF45[15];
    GRF45_16_buffer[clk] = GRF45[16];
    GRF45_17_buffer[clk] = GRF45[17];
    GRF45_18_buffer[clk] = GRF45[18];
    GRF45_19_buffer[clk] = GRF45[19];
    GRF45_20_buffer[clk] = GRF45[20];
    GRF45_21_buffer[clk] = GRF45[21];
    GRF45_22_buffer[clk] = GRF45[22];
    GRF45_23_buffer[clk] = GRF45[23];
    GRF45_24_buffer[clk] = GRF45[24];
    GRF45_25_buffer[clk] = GRF45[25];
    GRF45_26_buffer[clk] = GRF45[26];
    GRF45_27_buffer[clk] = GRF45[27];
    GRF45_28_buffer[clk] = GRF45[28];
    GRF45_29_buffer[clk] = GRF45[29];
    GRF45_30_buffer[clk] = GRF45[30];
    GRF45_31_buffer[clk] = GRF45[31];
    GRF46_0_buffer[clk] = GRF46[0];
    GRF46_1_buffer[clk] = GRF46[1];
    GRF46_2_buffer[clk] = GRF46[2];
    GRF46_3_buffer[clk] = GRF46[3];
    GRF46_4_buffer[clk] = GRF46[4];
    GRF46_5_buffer[clk] = GRF46[5];
    GRF46_6_buffer[clk] = GRF46[6];
    GRF46_7_buffer[clk] = GRF46[7];
    GRF46_8_buffer[clk] = GRF46[8];
    GRF46_9_buffer[clk] = GRF46[9];
    GRF46_10_buffer[clk] = GRF46[10];
    GRF46_11_buffer[clk] = GRF46[11];
    GRF46_12_buffer[clk] = GRF46[12];
    GRF46_13_buffer[clk] = GRF46[13];
    GRF46_14_buffer[clk] = GRF46[14];
    GRF46_15_buffer[clk] = GRF46[15];
    GRF46_16_buffer[clk] = GRF46[16];
    GRF46_17_buffer[clk] = GRF46[17];
    GRF46_18_buffer[clk] = GRF46[18];
    GRF46_19_buffer[clk] = GRF46[19];
    GRF46_20_buffer[clk] = GRF46[20];
    GRF46_21_buffer[clk] = GRF46[21];
    GRF46_22_buffer[clk] = GRF46[22];
    GRF46_23_buffer[clk] = GRF46[23];
    GRF46_24_buffer[clk] = GRF46[24];
    GRF46_25_buffer[clk] = GRF46[25];
    GRF46_26_buffer[clk] = GRF46[26];
    GRF46_27_buffer[clk] = GRF46[27];
    GRF46_28_buffer[clk] = GRF46[28];
    GRF46_29_buffer[clk] = GRF46[29];
    GRF46_30_buffer[clk] = GRF46[30];
    GRF46_31_buffer[clk] = GRF46[31];
    GRF47_0_buffer[clk] = GRF47[0];
    GRF47_1_buffer[clk] = GRF47[1];
    GRF47_2_buffer[clk] = GRF47[2];
    GRF47_3_buffer[clk] = GRF47[3];
    GRF47_4_buffer[clk] = GRF47[4];
    GRF47_5_buffer[clk] = GRF47[5];
    GRF47_6_buffer[clk] = GRF47[6];
    GRF47_7_buffer[clk] = GRF47[7];
    GRF47_8_buffer[clk] = GRF47[8];
    GRF47_9_buffer[clk] = GRF47[9];
    GRF47_10_buffer[clk] = GRF47[10];
    GRF47_11_buffer[clk] = GRF47[11];
    GRF47_12_buffer[clk] = GRF47[12];
    GRF47_13_buffer[clk] = GRF47[13];
    GRF47_14_buffer[clk] = GRF47[14];
    GRF47_15_buffer[clk] = GRF47[15];
    GRF47_16_buffer[clk] = GRF47[16];
    GRF47_17_buffer[clk] = GRF47[17];
    GRF47_18_buffer[clk] = GRF47[18];
    GRF47_19_buffer[clk] = GRF47[19];
    GRF47_20_buffer[clk] = GRF47[20];
    GRF47_21_buffer[clk] = GRF47[21];
    GRF47_22_buffer[clk] = GRF47[22];
    GRF47_23_buffer[clk] = GRF47[23];
    GRF47_24_buffer[clk] = GRF47[24];
    GRF47_25_buffer[clk] = GRF47[25];
    GRF47_26_buffer[clk] = GRF47[26];
    GRF47_27_buffer[clk] = GRF47[27];
    GRF47_28_buffer[clk] = GRF47[28];
    GRF47_29_buffer[clk] = GRF47[29];
    GRF47_30_buffer[clk] = GRF47[30];
    GRF47_31_buffer[clk] = GRF47[31];
    GRF48_0_buffer[clk] = GRF48[0];
    GRF48_1_buffer[clk] = GRF48[1];
    GRF48_2_buffer[clk] = GRF48[2];
    GRF48_3_buffer[clk] = GRF48[3];
    GRF48_4_buffer[clk] = GRF48[4];
    GRF48_5_buffer[clk] = GRF48[5];
    GRF48_6_buffer[clk] = GRF48[6];
    GRF48_7_buffer[clk] = GRF48[7];
    GRF48_8_buffer[clk] = GRF48[8];
    GRF48_9_buffer[clk] = GRF48[9];
    GRF48_10_buffer[clk] = GRF48[10];
    GRF48_11_buffer[clk] = GRF48[11];
    GRF48_12_buffer[clk] = GRF48[12];
    GRF48_13_buffer[clk] = GRF48[13];
    GRF48_14_buffer[clk] = GRF48[14];
    GRF48_15_buffer[clk] = GRF48[15];
    GRF48_16_buffer[clk] = GRF48[16];
    GRF48_17_buffer[clk] = GRF48[17];
    GRF48_18_buffer[clk] = GRF48[18];
    GRF48_19_buffer[clk] = GRF48[19];
    GRF48_20_buffer[clk] = GRF48[20];
    GRF48_21_buffer[clk] = GRF48[21];
    GRF48_22_buffer[clk] = GRF48[22];
    GRF48_23_buffer[clk] = GRF48[23];
    GRF48_24_buffer[clk] = GRF48[24];
    GRF48_25_buffer[clk] = GRF48[25];
    GRF48_26_buffer[clk] = GRF48[26];
    GRF48_27_buffer[clk] = GRF48[27];
    GRF48_28_buffer[clk] = GRF48[28];
    GRF48_29_buffer[clk] = GRF48[29];
    GRF48_30_buffer[clk] = GRF48[30];
    GRF48_31_buffer[clk] = GRF48[31];
    GRF49_0_buffer[clk] = GRF49[0];
    GRF49_1_buffer[clk] = GRF49[1];
    GRF49_2_buffer[clk] = GRF49[2];
    GRF49_3_buffer[clk] = GRF49[3];
    GRF49_4_buffer[clk] = GRF49[4];
    GRF49_5_buffer[clk] = GRF49[5];
    GRF49_6_buffer[clk] = GRF49[6];
    GRF49_7_buffer[clk] = GRF49[7];
    GRF49_8_buffer[clk] = GRF49[8];
    GRF49_9_buffer[clk] = GRF49[9];
    GRF49_10_buffer[clk] = GRF49[10];
    GRF49_11_buffer[clk] = GRF49[11];
    GRF49_12_buffer[clk] = GRF49[12];
    GRF49_13_buffer[clk] = GRF49[13];
    GRF49_14_buffer[clk] = GRF49[14];
    GRF49_15_buffer[clk] = GRF49[15];
    GRF49_16_buffer[clk] = GRF49[16];
    GRF49_17_buffer[clk] = GRF49[17];
    GRF49_18_buffer[clk] = GRF49[18];
    GRF49_19_buffer[clk] = GRF49[19];
    GRF49_20_buffer[clk] = GRF49[20];
    GRF49_21_buffer[clk] = GRF49[21];
    GRF49_22_buffer[clk] = GRF49[22];
    GRF49_23_buffer[clk] = GRF49[23];
    GRF49_24_buffer[clk] = GRF49[24];
    GRF49_25_buffer[clk] = GRF49[25];
    GRF49_26_buffer[clk] = GRF49[26];
    GRF49_27_buffer[clk] = GRF49[27];
    GRF49_28_buffer[clk] = GRF49[28];
    GRF49_29_buffer[clk] = GRF49[29];
    GRF49_30_buffer[clk] = GRF49[30];
    GRF49_31_buffer[clk] = GRF49[31];
    GRF50_0_buffer[clk] = GRF50[0];
    GRF50_1_buffer[clk] = GRF50[1];
    GRF50_2_buffer[clk] = GRF50[2];
    GRF50_3_buffer[clk] = GRF50[3];
    GRF50_4_buffer[clk] = GRF50[4];
    GRF50_5_buffer[clk] = GRF50[5];
    GRF50_6_buffer[clk] = GRF50[6];
    GRF50_7_buffer[clk] = GRF50[7];
    GRF50_8_buffer[clk] = GRF50[8];
    GRF50_9_buffer[clk] = GRF50[9];
    GRF50_10_buffer[clk] = GRF50[10];
    GRF50_11_buffer[clk] = GRF50[11];
    GRF50_12_buffer[clk] = GRF50[12];
    GRF50_13_buffer[clk] = GRF50[13];
    GRF50_14_buffer[clk] = GRF50[14];
    GRF50_15_buffer[clk] = GRF50[15];
    GRF50_16_buffer[clk] = GRF50[16];
    GRF50_17_buffer[clk] = GRF50[17];
    GRF50_18_buffer[clk] = GRF50[18];
    GRF50_19_buffer[clk] = GRF50[19];
    GRF50_20_buffer[clk] = GRF50[20];
    GRF50_21_buffer[clk] = GRF50[21];
    GRF50_22_buffer[clk] = GRF50[22];
    GRF50_23_buffer[clk] = GRF50[23];
    GRF50_24_buffer[clk] = GRF50[24];
    GRF50_25_buffer[clk] = GRF50[25];
    GRF50_26_buffer[clk] = GRF50[26];
    GRF50_27_buffer[clk] = GRF50[27];
    GRF50_28_buffer[clk] = GRF50[28];
    GRF50_29_buffer[clk] = GRF50[29];
    GRF50_30_buffer[clk] = GRF50[30];
    GRF50_31_buffer[clk] = GRF50[31];
    GRF51_0_buffer[clk] = GRF51[0];
    GRF51_1_buffer[clk] = GRF51[1];
    GRF51_2_buffer[clk] = GRF51[2];
    GRF51_3_buffer[clk] = GRF51[3];
    GRF51_4_buffer[clk] = GRF51[4];
    GRF51_5_buffer[clk] = GRF51[5];
    GRF51_6_buffer[clk] = GRF51[6];
    GRF51_7_buffer[clk] = GRF51[7];
    GRF51_8_buffer[clk] = GRF51[8];
    GRF51_9_buffer[clk] = GRF51[9];
    GRF51_10_buffer[clk] = GRF51[10];
    GRF51_11_buffer[clk] = GRF51[11];
    GRF51_12_buffer[clk] = GRF51[12];
    GRF51_13_buffer[clk] = GRF51[13];
    GRF51_14_buffer[clk] = GRF51[14];
    GRF51_15_buffer[clk] = GRF51[15];
    GRF51_16_buffer[clk] = GRF51[16];
    GRF51_17_buffer[clk] = GRF51[17];
    GRF51_18_buffer[clk] = GRF51[18];
    GRF51_19_buffer[clk] = GRF51[19];
    GRF51_20_buffer[clk] = GRF51[20];
    GRF51_21_buffer[clk] = GRF51[21];
    GRF51_22_buffer[clk] = GRF51[22];
    GRF51_23_buffer[clk] = GRF51[23];
    GRF51_24_buffer[clk] = GRF51[24];
    GRF51_25_buffer[clk] = GRF51[25];
    GRF51_26_buffer[clk] = GRF51[26];
    GRF51_27_buffer[clk] = GRF51[27];
    GRF51_28_buffer[clk] = GRF51[28];
    GRF51_29_buffer[clk] = GRF51[29];
    GRF51_30_buffer[clk] = GRF51[30];
    GRF51_31_buffer[clk] = GRF51[31];
    GRF52_0_buffer[clk] = GRF52[0];
    GRF52_1_buffer[clk] = GRF52[1];
    GRF52_2_buffer[clk] = GRF52[2];
    GRF52_3_buffer[clk] = GRF52[3];
    GRF52_4_buffer[clk] = GRF52[4];
    GRF52_5_buffer[clk] = GRF52[5];
    GRF52_6_buffer[clk] = GRF52[6];
    GRF52_7_buffer[clk] = GRF52[7];
    GRF52_8_buffer[clk] = GRF52[8];
    GRF52_9_buffer[clk] = GRF52[9];
    GRF52_10_buffer[clk] = GRF52[10];
    GRF52_11_buffer[clk] = GRF52[11];
    GRF52_12_buffer[clk] = GRF52[12];
    GRF52_13_buffer[clk] = GRF52[13];
    GRF52_14_buffer[clk] = GRF52[14];
    GRF52_15_buffer[clk] = GRF52[15];
    GRF52_16_buffer[clk] = GRF52[16];
    GRF52_17_buffer[clk] = GRF52[17];
    GRF52_18_buffer[clk] = GRF52[18];
    GRF52_19_buffer[clk] = GRF52[19];
    GRF52_20_buffer[clk] = GRF52[20];
    GRF52_21_buffer[clk] = GRF52[21];
    GRF52_22_buffer[clk] = GRF52[22];
    GRF52_23_buffer[clk] = GRF52[23];
    GRF52_24_buffer[clk] = GRF52[24];
    GRF52_25_buffer[clk] = GRF52[25];
    GRF52_26_buffer[clk] = GRF52[26];
    GRF52_27_buffer[clk] = GRF52[27];
    GRF52_28_buffer[clk] = GRF52[28];
    GRF52_29_buffer[clk] = GRF52[29];
    GRF52_30_buffer[clk] = GRF52[30];
    GRF52_31_buffer[clk] = GRF52[31];
    GRF53_0_buffer[clk] = GRF53[0];
    GRF53_1_buffer[clk] = GRF53[1];
    GRF53_2_buffer[clk] = GRF53[2];
    GRF53_3_buffer[clk] = GRF53[3];
    GRF53_4_buffer[clk] = GRF53[4];
    GRF53_5_buffer[clk] = GRF53[5];
    GRF53_6_buffer[clk] = GRF53[6];
    GRF53_7_buffer[clk] = GRF53[7];
    GRF53_8_buffer[clk] = GRF53[8];
    GRF53_9_buffer[clk] = GRF53[9];
    GRF53_10_buffer[clk] = GRF53[10];
    GRF53_11_buffer[clk] = GRF53[11];
    GRF53_12_buffer[clk] = GRF53[12];
    GRF53_13_buffer[clk] = GRF53[13];
    GRF53_14_buffer[clk] = GRF53[14];
    GRF53_15_buffer[clk] = GRF53[15];
    GRF53_16_buffer[clk] = GRF53[16];
    GRF53_17_buffer[clk] = GRF53[17];
    GRF53_18_buffer[clk] = GRF53[18];
    GRF53_19_buffer[clk] = GRF53[19];
    GRF53_20_buffer[clk] = GRF53[20];
    GRF53_21_buffer[clk] = GRF53[21];
    GRF53_22_buffer[clk] = GRF53[22];
    GRF53_23_buffer[clk] = GRF53[23];
    GRF53_24_buffer[clk] = GRF53[24];
    GRF53_25_buffer[clk] = GRF53[25];
    GRF53_26_buffer[clk] = GRF53[26];
    GRF53_27_buffer[clk] = GRF53[27];
    GRF53_28_buffer[clk] = GRF53[28];
    GRF53_29_buffer[clk] = GRF53[29];
    GRF53_30_buffer[clk] = GRF53[30];
    GRF53_31_buffer[clk] = GRF53[31];
    GRF54_0_buffer[clk] = GRF54[0];
    GRF54_1_buffer[clk] = GRF54[1];
    GRF54_2_buffer[clk] = GRF54[2];
    GRF54_3_buffer[clk] = GRF54[3];
    GRF54_4_buffer[clk] = GRF54[4];
    GRF54_5_buffer[clk] = GRF54[5];
    GRF54_6_buffer[clk] = GRF54[6];
    GRF54_7_buffer[clk] = GRF54[7];
    GRF54_8_buffer[clk] = GRF54[8];
    GRF54_9_buffer[clk] = GRF54[9];
    GRF54_10_buffer[clk] = GRF54[10];
    GRF54_11_buffer[clk] = GRF54[11];
    GRF54_12_buffer[clk] = GRF54[12];
    GRF54_13_buffer[clk] = GRF54[13];
    GRF54_14_buffer[clk] = GRF54[14];
    GRF54_15_buffer[clk] = GRF54[15];
    GRF54_16_buffer[clk] = GRF54[16];
    GRF54_17_buffer[clk] = GRF54[17];
    GRF54_18_buffer[clk] = GRF54[18];
    GRF54_19_buffer[clk] = GRF54[19];
    GRF54_20_buffer[clk] = GRF54[20];
    GRF54_21_buffer[clk] = GRF54[21];
    GRF54_22_buffer[clk] = GRF54[22];
    GRF54_23_buffer[clk] = GRF54[23];
    GRF54_24_buffer[clk] = GRF54[24];
    GRF54_25_buffer[clk] = GRF54[25];
    GRF54_26_buffer[clk] = GRF54[26];
    GRF54_27_buffer[clk] = GRF54[27];
    GRF54_28_buffer[clk] = GRF54[28];
    GRF54_29_buffer[clk] = GRF54[29];
    GRF54_30_buffer[clk] = GRF54[30];
    GRF54_31_buffer[clk] = GRF54[31];
    GRF55_0_buffer[clk] = GRF55[0];
    GRF55_1_buffer[clk] = GRF55[1];
    GRF55_2_buffer[clk] = GRF55[2];
    GRF55_3_buffer[clk] = GRF55[3];
    GRF55_4_buffer[clk] = GRF55[4];
    GRF55_5_buffer[clk] = GRF55[5];
    GRF55_6_buffer[clk] = GRF55[6];
    GRF55_7_buffer[clk] = GRF55[7];
    GRF55_8_buffer[clk] = GRF55[8];
    GRF55_9_buffer[clk] = GRF55[9];
    GRF55_10_buffer[clk] = GRF55[10];
    GRF55_11_buffer[clk] = GRF55[11];
    GRF55_12_buffer[clk] = GRF55[12];
    GRF55_13_buffer[clk] = GRF55[13];
    GRF55_14_buffer[clk] = GRF55[14];
    GRF55_15_buffer[clk] = GRF55[15];
    GRF55_16_buffer[clk] = GRF55[16];
    GRF55_17_buffer[clk] = GRF55[17];
    GRF55_18_buffer[clk] = GRF55[18];
    GRF55_19_buffer[clk] = GRF55[19];
    GRF55_20_buffer[clk] = GRF55[20];
    GRF55_21_buffer[clk] = GRF55[21];
    GRF55_22_buffer[clk] = GRF55[22];
    GRF55_23_buffer[clk] = GRF55[23];
    GRF55_24_buffer[clk] = GRF55[24];
    GRF55_25_buffer[clk] = GRF55[25];
    GRF55_26_buffer[clk] = GRF55[26];
    GRF55_27_buffer[clk] = GRF55[27];
    GRF55_28_buffer[clk] = GRF55[28];
    GRF55_29_buffer[clk] = GRF55[29];
    GRF55_30_buffer[clk] = GRF55[30];
    GRF55_31_buffer[clk] = GRF55[31];
    GRF56_0_buffer[clk] = GRF56[0];
    GRF56_1_buffer[clk] = GRF56[1];
    GRF56_2_buffer[clk] = GRF56[2];
    GRF56_3_buffer[clk] = GRF56[3];
    GRF56_4_buffer[clk] = GRF56[4];
    GRF56_5_buffer[clk] = GRF56[5];
    GRF56_6_buffer[clk] = GRF56[6];
    GRF56_7_buffer[clk] = GRF56[7];
    GRF56_8_buffer[clk] = GRF56[8];
    GRF56_9_buffer[clk] = GRF56[9];
    GRF56_10_buffer[clk] = GRF56[10];
    GRF56_11_buffer[clk] = GRF56[11];
    GRF56_12_buffer[clk] = GRF56[12];
    GRF56_13_buffer[clk] = GRF56[13];
    GRF56_14_buffer[clk] = GRF56[14];
    GRF56_15_buffer[clk] = GRF56[15];
    GRF56_16_buffer[clk] = GRF56[16];
    GRF56_17_buffer[clk] = GRF56[17];
    GRF56_18_buffer[clk] = GRF56[18];
    GRF56_19_buffer[clk] = GRF56[19];
    GRF56_20_buffer[clk] = GRF56[20];
    GRF56_21_buffer[clk] = GRF56[21];
    GRF56_22_buffer[clk] = GRF56[22];
    GRF56_23_buffer[clk] = GRF56[23];
    GRF56_24_buffer[clk] = GRF56[24];
    GRF56_25_buffer[clk] = GRF56[25];
    GRF56_26_buffer[clk] = GRF56[26];
    GRF56_27_buffer[clk] = GRF56[27];
    GRF56_28_buffer[clk] = GRF56[28];
    GRF56_29_buffer[clk] = GRF56[29];
    GRF56_30_buffer[clk] = GRF56[30];
    GRF56_31_buffer[clk] = GRF56[31];
    GRF57_0_buffer[clk] = GRF57[0];
    GRF57_1_buffer[clk] = GRF57[1];
    GRF57_2_buffer[clk] = GRF57[2];
    GRF57_3_buffer[clk] = GRF57[3];
    GRF57_4_buffer[clk] = GRF57[4];
    GRF57_5_buffer[clk] = GRF57[5];
    GRF57_6_buffer[clk] = GRF57[6];
    GRF57_7_buffer[clk] = GRF57[7];
    GRF57_8_buffer[clk] = GRF57[8];
    GRF57_9_buffer[clk] = GRF57[9];
    GRF57_10_buffer[clk] = GRF57[10];
    GRF57_11_buffer[clk] = GRF57[11];
    GRF57_12_buffer[clk] = GRF57[12];
    GRF57_13_buffer[clk] = GRF57[13];
    GRF57_14_buffer[clk] = GRF57[14];
    GRF57_15_buffer[clk] = GRF57[15];
    GRF57_16_buffer[clk] = GRF57[16];
    GRF57_17_buffer[clk] = GRF57[17];
    GRF57_18_buffer[clk] = GRF57[18];
    GRF57_19_buffer[clk] = GRF57[19];
    GRF57_20_buffer[clk] = GRF57[20];
    GRF57_21_buffer[clk] = GRF57[21];
    GRF57_22_buffer[clk] = GRF57[22];
    GRF57_23_buffer[clk] = GRF57[23];
    GRF57_24_buffer[clk] = GRF57[24];
    GRF57_25_buffer[clk] = GRF57[25];
    GRF57_26_buffer[clk] = GRF57[26];
    GRF57_27_buffer[clk] = GRF57[27];
    GRF57_28_buffer[clk] = GRF57[28];
    GRF57_29_buffer[clk] = GRF57[29];
    GRF57_30_buffer[clk] = GRF57[30];
    GRF57_31_buffer[clk] = GRF57[31];
    GRF58_0_buffer[clk] = GRF58[0];
    GRF58_1_buffer[clk] = GRF58[1];
    GRF58_2_buffer[clk] = GRF58[2];
    GRF58_3_buffer[clk] = GRF58[3];
    GRF58_4_buffer[clk] = GRF58[4];
    GRF58_5_buffer[clk] = GRF58[5];
    GRF58_6_buffer[clk] = GRF58[6];
    GRF58_7_buffer[clk] = GRF58[7];
    GRF58_8_buffer[clk] = GRF58[8];
    GRF58_9_buffer[clk] = GRF58[9];
    GRF58_10_buffer[clk] = GRF58[10];
    GRF58_11_buffer[clk] = GRF58[11];
    GRF58_12_buffer[clk] = GRF58[12];
    GRF58_13_buffer[clk] = GRF58[13];
    GRF58_14_buffer[clk] = GRF58[14];
    GRF58_15_buffer[clk] = GRF58[15];
    GRF58_16_buffer[clk] = GRF58[16];
    GRF58_17_buffer[clk] = GRF58[17];
    GRF58_18_buffer[clk] = GRF58[18];
    GRF58_19_buffer[clk] = GRF58[19];
    GRF58_20_buffer[clk] = GRF58[20];
    GRF58_21_buffer[clk] = GRF58[21];
    GRF58_22_buffer[clk] = GRF58[22];
    GRF58_23_buffer[clk] = GRF58[23];
    GRF58_24_buffer[clk] = GRF58[24];
    GRF58_25_buffer[clk] = GRF58[25];
    GRF58_26_buffer[clk] = GRF58[26];
    GRF58_27_buffer[clk] = GRF58[27];
    GRF58_28_buffer[clk] = GRF58[28];
    GRF58_29_buffer[clk] = GRF58[29];
    GRF58_30_buffer[clk] = GRF58[30];
    GRF58_31_buffer[clk] = GRF58[31];
    GRF59_0_buffer[clk] = GRF59[0];
    GRF59_1_buffer[clk] = GRF59[1];
    GRF59_2_buffer[clk] = GRF59[2];
    GRF59_3_buffer[clk] = GRF59[3];
    GRF59_4_buffer[clk] = GRF59[4];
    GRF59_5_buffer[clk] = GRF59[5];
    GRF59_6_buffer[clk] = GRF59[6];
    GRF59_7_buffer[clk] = GRF59[7];
    GRF59_8_buffer[clk] = GRF59[8];
    GRF59_9_buffer[clk] = GRF59[9];
    GRF59_10_buffer[clk] = GRF59[10];
    GRF59_11_buffer[clk] = GRF59[11];
    GRF59_12_buffer[clk] = GRF59[12];
    GRF59_13_buffer[clk] = GRF59[13];
    GRF59_14_buffer[clk] = GRF59[14];
    GRF59_15_buffer[clk] = GRF59[15];
    GRF59_16_buffer[clk] = GRF59[16];
    GRF59_17_buffer[clk] = GRF59[17];
    GRF59_18_buffer[clk] = GRF59[18];
    GRF59_19_buffer[clk] = GRF59[19];
    GRF59_20_buffer[clk] = GRF59[20];
    GRF59_21_buffer[clk] = GRF59[21];
    GRF59_22_buffer[clk] = GRF59[22];
    GRF59_23_buffer[clk] = GRF59[23];
    GRF59_24_buffer[clk] = GRF59[24];
    GRF59_25_buffer[clk] = GRF59[25];
    GRF59_26_buffer[clk] = GRF59[26];
    GRF59_27_buffer[clk] = GRF59[27];
    GRF59_28_buffer[clk] = GRF59[28];
    GRF59_29_buffer[clk] = GRF59[29];
    GRF59_30_buffer[clk] = GRF59[30];
    GRF59_31_buffer[clk] = GRF59[31];
    GRF60_0_buffer[clk] = GRF60[0];
    GRF60_1_buffer[clk] = GRF60[1];
    GRF60_2_buffer[clk] = GRF60[2];
    GRF60_3_buffer[clk] = GRF60[3];
    GRF60_4_buffer[clk] = GRF60[4];
    GRF60_5_buffer[clk] = GRF60[5];
    GRF60_6_buffer[clk] = GRF60[6];
    GRF60_7_buffer[clk] = GRF60[7];
    GRF60_8_buffer[clk] = GRF60[8];
    GRF60_9_buffer[clk] = GRF60[9];
    GRF60_10_buffer[clk] = GRF60[10];
    GRF60_11_buffer[clk] = GRF60[11];
    GRF60_12_buffer[clk] = GRF60[12];
    GRF60_13_buffer[clk] = GRF60[13];
    GRF60_14_buffer[clk] = GRF60[14];
    GRF60_15_buffer[clk] = GRF60[15];
    GRF60_16_buffer[clk] = GRF60[16];
    GRF60_17_buffer[clk] = GRF60[17];
    GRF60_18_buffer[clk] = GRF60[18];
    GRF60_19_buffer[clk] = GRF60[19];
    GRF60_20_buffer[clk] = GRF60[20];
    GRF60_21_buffer[clk] = GRF60[21];
    GRF60_22_buffer[clk] = GRF60[22];
    GRF60_23_buffer[clk] = GRF60[23];
    GRF60_24_buffer[clk] = GRF60[24];
    GRF60_25_buffer[clk] = GRF60[25];
    GRF60_26_buffer[clk] = GRF60[26];
    GRF60_27_buffer[clk] = GRF60[27];
    GRF60_28_buffer[clk] = GRF60[28];
    GRF60_29_buffer[clk] = GRF60[29];
    GRF60_30_buffer[clk] = GRF60[30];
    GRF60_31_buffer[clk] = GRF60[31];
    GRF61_0_buffer[clk] = GRF61[0];
    GRF61_1_buffer[clk] = GRF61[1];
    GRF61_2_buffer[clk] = GRF61[2];
    GRF61_3_buffer[clk] = GRF61[3];
    GRF61_4_buffer[clk] = GRF61[4];
    GRF61_5_buffer[clk] = GRF61[5];
    GRF61_6_buffer[clk] = GRF61[6];
    GRF61_7_buffer[clk] = GRF61[7];
    GRF61_8_buffer[clk] = GRF61[8];
    GRF61_9_buffer[clk] = GRF61[9];
    GRF61_10_buffer[clk] = GRF61[10];
    GRF61_11_buffer[clk] = GRF61[11];
    GRF61_12_buffer[clk] = GRF61[12];
    GRF61_13_buffer[clk] = GRF61[13];
    GRF61_14_buffer[clk] = GRF61[14];
    GRF61_15_buffer[clk] = GRF61[15];
    GRF61_16_buffer[clk] = GRF61[16];
    GRF61_17_buffer[clk] = GRF61[17];
    GRF61_18_buffer[clk] = GRF61[18];
    GRF61_19_buffer[clk] = GRF61[19];
    GRF61_20_buffer[clk] = GRF61[20];
    GRF61_21_buffer[clk] = GRF61[21];
    GRF61_22_buffer[clk] = GRF61[22];
    GRF61_23_buffer[clk] = GRF61[23];
    GRF61_24_buffer[clk] = GRF61[24];
    GRF61_25_buffer[clk] = GRF61[25];
    GRF61_26_buffer[clk] = GRF61[26];
    GRF61_27_buffer[clk] = GRF61[27];
    GRF61_28_buffer[clk] = GRF61[28];
    GRF61_29_buffer[clk] = GRF61[29];
    GRF61_30_buffer[clk] = GRF61[30];
    GRF61_31_buffer[clk] = GRF61[31];
    GRF62_0_buffer[clk] = GRF62[0];
    GRF62_1_buffer[clk] = GRF62[1];
    GRF62_2_buffer[clk] = GRF62[2];
    GRF62_3_buffer[clk] = GRF62[3];
    GRF62_4_buffer[clk] = GRF62[4];
    GRF62_5_buffer[clk] = GRF62[5];
    GRF62_6_buffer[clk] = GRF62[6];
    GRF62_7_buffer[clk] = GRF62[7];
    GRF62_8_buffer[clk] = GRF62[8];
    GRF62_9_buffer[clk] = GRF62[9];
    GRF62_10_buffer[clk] = GRF62[10];
    GRF62_11_buffer[clk] = GRF62[11];
    GRF62_12_buffer[clk] = GRF62[12];
    GRF62_13_buffer[clk] = GRF62[13];
    GRF62_14_buffer[clk] = GRF62[14];
    GRF62_15_buffer[clk] = GRF62[15];
    GRF62_16_buffer[clk] = GRF62[16];
    GRF62_17_buffer[clk] = GRF62[17];
    GRF62_18_buffer[clk] = GRF62[18];
    GRF62_19_buffer[clk] = GRF62[19];
    GRF62_20_buffer[clk] = GRF62[20];
    GRF62_21_buffer[clk] = GRF62[21];
    GRF62_22_buffer[clk] = GRF62[22];
    GRF62_23_buffer[clk] = GRF62[23];
    GRF62_24_buffer[clk] = GRF62[24];
    GRF62_25_buffer[clk] = GRF62[25];
    GRF62_26_buffer[clk] = GRF62[26];
    GRF62_27_buffer[clk] = GRF62[27];
    GRF62_28_buffer[clk] = GRF62[28];
    GRF62_29_buffer[clk] = GRF62[29];
    GRF62_30_buffer[clk] = GRF62[30];
    GRF62_31_buffer[clk] = GRF62[31];
    GRF63_0_buffer[clk] = GRF63[0];
    GRF63_1_buffer[clk] = GRF63[1];
    GRF63_2_buffer[clk] = GRF63[2];
    GRF63_3_buffer[clk] = GRF63[3];
    GRF63_4_buffer[clk] = GRF63[4];
    GRF63_5_buffer[clk] = GRF63[5];
    GRF63_6_buffer[clk] = GRF63[6];
    GRF63_7_buffer[clk] = GRF63[7];
    GRF63_8_buffer[clk] = GRF63[8];
    GRF63_9_buffer[clk] = GRF63[9];
    GRF63_10_buffer[clk] = GRF63[10];
    GRF63_11_buffer[clk] = GRF63[11];
    GRF63_12_buffer[clk] = GRF63[12];
    GRF63_13_buffer[clk] = GRF63[13];
    GRF63_14_buffer[clk] = GRF63[14];
    GRF63_15_buffer[clk] = GRF63[15];
    GRF63_16_buffer[clk] = GRF63[16];
    GRF63_17_buffer[clk] = GRF63[17];
    GRF63_18_buffer[clk] = GRF63[18];
    GRF63_19_buffer[clk] = GRF63[19];
    GRF63_20_buffer[clk] = GRF63[20];
    GRF63_21_buffer[clk] = GRF63[21];
    GRF63_22_buffer[clk] = GRF63[22];
    GRF63_23_buffer[clk] = GRF63[23];
    GRF63_24_buffer[clk] = GRF63[24];
    GRF63_25_buffer[clk] = GRF63[25];
    GRF63_26_buffer[clk] = GRF63[26];
    GRF63_27_buffer[clk] = GRF63[27];
    GRF63_28_buffer[clk] = GRF63[28];
    GRF63_29_buffer[clk] = GRF63[29];
    GRF63_30_buffer[clk] = GRF63[30];
    GRF63_31_buffer[clk] = GRF63[31];
  end


  // generate warp signal 
  always_comb begin
    if ((GRF0_0_buffer[clk] != GRF0_0_buffer[!clk]) ||(GRF0_1_buffer[clk] != GRF0_1_buffer[!clk]) ||(GRF0_2_buffer[clk] != GRF0_2_buffer[!clk]) ||(GRF0_3_buffer[clk] != GRF0_3_buffer[!clk]) ||(GRF0_4_buffer[clk] != GRF0_4_buffer[!clk]) ||(GRF0_5_buffer[clk] != GRF0_5_buffer[!clk]) ||(GRF0_6_buffer[clk] != GRF0_6_buffer[!clk]) ||(GRF0_7_buffer[clk] != GRF0_7_buffer[!clk]) ||(GRF0_8_buffer[clk] != GRF0_8_buffer[!clk]) ||(GRF0_9_buffer[clk] != GRF0_9_buffer[!clk]) ||(GRF0_10_buffer[clk] != GRF0_10_buffer[!clk]) ||(GRF0_11_buffer[clk] != GRF0_11_buffer[!clk]) ||(GRF0_12_buffer[clk] != GRF0_12_buffer[!clk]) ||(GRF0_13_buffer[clk] != GRF0_13_buffer[!clk]) ||(GRF0_14_buffer[clk] != GRF0_14_buffer[!clk]) ||(GRF0_15_buffer[clk] != GRF0_15_buffer[!clk]) ||(GRF0_16_buffer[clk] != GRF0_16_buffer[!clk]) ||(GRF0_17_buffer[clk] != GRF0_17_buffer[!clk]) ||(GRF0_18_buffer[clk] != GRF0_18_buffer[!clk]) ||(GRF0_19_buffer[clk] != GRF0_19_buffer[!clk]) ||(GRF0_20_buffer[clk] != GRF0_20_buffer[!clk]) ||(GRF0_21_buffer[clk] != GRF0_21_buffer[!clk]) ||(GRF0_22_buffer[clk] != GRF0_22_buffer[!clk]) ||(GRF0_23_buffer[clk] != GRF0_23_buffer[!clk]) ||(GRF0_24_buffer[clk] != GRF0_24_buffer[!clk]) ||(GRF0_25_buffer[clk] != GRF0_25_buffer[!clk]) ||(GRF0_26_buffer[clk] != GRF0_26_buffer[!clk]) ||(GRF0_27_buffer[clk] != GRF0_27_buffer[!clk]) ||(GRF0_28_buffer[clk] != GRF0_28_buffer[!clk]) ||(GRF0_29_buffer[clk] != GRF0_29_buffer[!clk]) ||(GRF0_30_buffer[clk] != GRF0_30_buffer[!clk]) ||(GRF0_31_buffer[clk] != GRF0_31_buffer[!clk]) ||(GRF8_0_buffer[clk] != GRF8_0_buffer[!clk]) ||(GRF8_1_buffer[clk] != GRF8_1_buffer[!clk]) ||(GRF8_2_buffer[clk] != GRF8_2_buffer[!clk]) ||(GRF8_3_buffer[clk] != GRF8_3_buffer[!clk]) ||(GRF8_4_buffer[clk] != GRF8_4_buffer[!clk]) ||(GRF8_5_buffer[clk] != GRF8_5_buffer[!clk]) ||(GRF8_6_buffer[clk] != GRF8_6_buffer[!clk]) ||(GRF8_7_buffer[clk] != GRF8_7_buffer[!clk]) ||(GRF8_8_buffer[clk] != GRF8_8_buffer[!clk]) ||(GRF8_9_buffer[clk] != GRF8_9_buffer[!clk]) ||(GRF8_10_buffer[clk] != GRF8_10_buffer[!clk]) ||(GRF8_11_buffer[clk] != GRF8_11_buffer[!clk]) ||(GRF8_12_buffer[clk] != GRF8_12_buffer[!clk]) ||(GRF8_13_buffer[clk] != GRF8_13_buffer[!clk]) ||(GRF8_14_buffer[clk] != GRF8_14_buffer[!clk]) ||(GRF8_15_buffer[clk] != GRF8_15_buffer[!clk]) ||(GRF8_16_buffer[clk] != GRF8_16_buffer[!clk]) ||(GRF8_17_buffer[clk] != GRF8_17_buffer[!clk]) ||(GRF8_18_buffer[clk] != GRF8_18_buffer[!clk]) ||(GRF8_19_buffer[clk] != GRF8_19_buffer[!clk]) ||(GRF8_20_buffer[clk] != GRF8_20_buffer[!clk]) ||(GRF8_21_buffer[clk] != GRF8_21_buffer[!clk]) ||(GRF8_22_buffer[clk] != GRF8_22_buffer[!clk]) ||(GRF8_23_buffer[clk] != GRF8_23_buffer[!clk]) ||(GRF8_24_buffer[clk] != GRF8_24_buffer[!clk]) ||(GRF8_25_buffer[clk] != GRF8_25_buffer[!clk]) ||(GRF8_26_buffer[clk] != GRF8_26_buffer[!clk]) ||(GRF8_27_buffer[clk] != GRF8_27_buffer[!clk]) ||(GRF8_28_buffer[clk] != GRF8_28_buffer[!clk]) ||(GRF8_29_buffer[clk] != GRF8_29_buffer[!clk]) ||(GRF8_30_buffer[clk] != GRF8_30_buffer[!clk]) ||(GRF8_31_buffer[clk] != GRF8_31_buffer[!clk]) ||(GRF16_0_buffer[clk] != GRF16_0_buffer[!clk]) ||(GRF16_1_buffer[clk] != GRF16_1_buffer[!clk]) ||(GRF16_2_buffer[clk] != GRF16_2_buffer[!clk]) ||(GRF16_3_buffer[clk] != GRF16_3_buffer[!clk]) ||(GRF16_4_buffer[clk] != GRF16_4_buffer[!clk]) ||(GRF16_5_buffer[clk] != GRF16_5_buffer[!clk]) ||(GRF16_6_buffer[clk] != GRF16_6_buffer[!clk]) ||(GRF16_7_buffer[clk] != GRF16_7_buffer[!clk]) ||(GRF16_8_buffer[clk] != GRF16_8_buffer[!clk]) ||(GRF16_9_buffer[clk] != GRF16_9_buffer[!clk]) ||(GRF16_10_buffer[clk] != GRF16_10_buffer[!clk]) ||(GRF16_11_buffer[clk] != GRF16_11_buffer[!clk]) ||(GRF16_12_buffer[clk] != GRF16_12_buffer[!clk]) ||(GRF16_13_buffer[clk] != GRF16_13_buffer[!clk]) ||(GRF16_14_buffer[clk] != GRF16_14_buffer[!clk]) ||(GRF16_15_buffer[clk] != GRF16_15_buffer[!clk]) ||(GRF16_16_buffer[clk] != GRF16_16_buffer[!clk]) ||(GRF16_17_buffer[clk] != GRF16_17_buffer[!clk]) ||(GRF16_18_buffer[clk] != GRF16_18_buffer[!clk]) ||(GRF16_19_buffer[clk] != GRF16_19_buffer[!clk]) ||(GRF16_20_buffer[clk] != GRF16_20_buffer[!clk]) ||(GRF16_21_buffer[clk] != GRF16_21_buffer[!clk]) ||(GRF16_22_buffer[clk] != GRF16_22_buffer[!clk]) ||(GRF16_23_buffer[clk] != GRF16_23_buffer[!clk]) ||(GRF16_24_buffer[clk] != GRF16_24_buffer[!clk]) ||(GRF16_25_buffer[clk] != GRF16_25_buffer[!clk]) ||(GRF16_26_buffer[clk] != GRF16_26_buffer[!clk]) ||(GRF16_27_buffer[clk] != GRF16_27_buffer[!clk]) ||(GRF16_28_buffer[clk] != GRF16_28_buffer[!clk]) ||(GRF16_29_buffer[clk] != GRF16_29_buffer[!clk]) ||(GRF16_30_buffer[clk] != GRF16_30_buffer[!clk]) ||(GRF16_31_buffer[clk] != GRF16_31_buffer[!clk]) ||(GRF24_0_buffer[clk] != GRF24_0_buffer[!clk]) ||(GRF24_1_buffer[clk] != GRF24_1_buffer[!clk]) ||(GRF24_2_buffer[clk] != GRF24_2_buffer[!clk]) ||(GRF24_3_buffer[clk] != GRF24_3_buffer[!clk]) ||(GRF24_4_buffer[clk] != GRF24_4_buffer[!clk]) ||(GRF24_5_buffer[clk] != GRF24_5_buffer[!clk]) ||(GRF24_6_buffer[clk] != GRF24_6_buffer[!clk]) ||(GRF24_7_buffer[clk] != GRF24_7_buffer[!clk]) ||(GRF24_8_buffer[clk] != GRF24_8_buffer[!clk]) ||(GRF24_9_buffer[clk] != GRF24_9_buffer[!clk]) ||(GRF24_10_buffer[clk] != GRF24_10_buffer[!clk]) ||(GRF24_11_buffer[clk] != GRF24_11_buffer[!clk]) ||(GRF24_12_buffer[clk] != GRF24_12_buffer[!clk]) ||(GRF24_13_buffer[clk] != GRF24_13_buffer[!clk]) ||(GRF24_14_buffer[clk] != GRF24_14_buffer[!clk]) ||(GRF24_15_buffer[clk] != GRF24_15_buffer[!clk]) ||(GRF24_16_buffer[clk] != GRF24_16_buffer[!clk]) ||(GRF24_17_buffer[clk] != GRF24_17_buffer[!clk]) ||(GRF24_18_buffer[clk] != GRF24_18_buffer[!clk]) ||(GRF24_19_buffer[clk] != GRF24_19_buffer[!clk]) ||(GRF24_20_buffer[clk] != GRF24_20_buffer[!clk]) ||(GRF24_21_buffer[clk] != GRF24_21_buffer[!clk]) ||(GRF24_22_buffer[clk] != GRF24_22_buffer[!clk]) ||(GRF24_23_buffer[clk] != GRF24_23_buffer[!clk]) ||(GRF24_24_buffer[clk] != GRF24_24_buffer[!clk]) ||(GRF24_25_buffer[clk] != GRF24_25_buffer[!clk]) ||(GRF24_26_buffer[clk] != GRF24_26_buffer[!clk]) ||(GRF24_27_buffer[clk] != GRF24_27_buffer[!clk]) ||(GRF24_28_buffer[clk] != GRF24_28_buffer[!clk]) ||(GRF24_29_buffer[clk] != GRF24_29_buffer[!clk]) ||(GRF24_30_buffer[clk] != GRF24_30_buffer[!clk]) ||(GRF24_31_buffer[clk] != GRF24_31_buffer[!clk]) ||(GRF32_0_buffer[clk] != GRF32_0_buffer[!clk]) ||(GRF32_1_buffer[clk] != GRF32_1_buffer[!clk]) ||(GRF32_2_buffer[clk] != GRF32_2_buffer[!clk]) ||(GRF32_3_buffer[clk] != GRF32_3_buffer[!clk]) ||(GRF32_4_buffer[clk] != GRF32_4_buffer[!clk]) ||(GRF32_5_buffer[clk] != GRF32_5_buffer[!clk]) ||(GRF32_6_buffer[clk] != GRF32_6_buffer[!clk]) ||(GRF32_7_buffer[clk] != GRF32_7_buffer[!clk]) ||(GRF32_8_buffer[clk] != GRF32_8_buffer[!clk]) ||(GRF32_9_buffer[clk] != GRF32_9_buffer[!clk]) ||(GRF32_10_buffer[clk] != GRF32_10_buffer[!clk]) ||(GRF32_11_buffer[clk] != GRF32_11_buffer[!clk]) ||(GRF32_12_buffer[clk] != GRF32_12_buffer[!clk]) ||(GRF32_13_buffer[clk] != GRF32_13_buffer[!clk]) ||(GRF32_14_buffer[clk] != GRF32_14_buffer[!clk]) ||(GRF32_15_buffer[clk] != GRF32_15_buffer[!clk]) ||(GRF32_16_buffer[clk] != GRF32_16_buffer[!clk]) ||(GRF32_17_buffer[clk] != GRF32_17_buffer[!clk]) ||(GRF32_18_buffer[clk] != GRF32_18_buffer[!clk]) ||(GRF32_19_buffer[clk] != GRF32_19_buffer[!clk]) ||(GRF32_20_buffer[clk] != GRF32_20_buffer[!clk]) ||(GRF32_21_buffer[clk] != GRF32_21_buffer[!clk]) ||(GRF32_22_buffer[clk] != GRF32_22_buffer[!clk]) ||(GRF32_23_buffer[clk] != GRF32_23_buffer[!clk]) ||(GRF32_24_buffer[clk] != GRF32_24_buffer[!clk]) ||(GRF32_25_buffer[clk] != GRF32_25_buffer[!clk]) ||(GRF32_26_buffer[clk] != GRF32_26_buffer[!clk]) ||(GRF32_27_buffer[clk] != GRF32_27_buffer[!clk]) ||(GRF32_28_buffer[clk] != GRF32_28_buffer[!clk]) ||(GRF32_29_buffer[clk] != GRF32_29_buffer[!clk]) ||(GRF32_30_buffer[clk] != GRF32_30_buffer[!clk]) ||(GRF32_31_buffer[clk] != GRF32_31_buffer[!clk]) ||(GRF40_0_buffer[clk] != GRF40_0_buffer[!clk]) ||(GRF40_1_buffer[clk] != GRF40_1_buffer[!clk]) ||(GRF40_2_buffer[clk] != GRF40_2_buffer[!clk]) ||(GRF40_3_buffer[clk] != GRF40_3_buffer[!clk]) ||(GRF40_4_buffer[clk] != GRF40_4_buffer[!clk]) ||(GRF40_5_buffer[clk] != GRF40_5_buffer[!clk]) ||(GRF40_6_buffer[clk] != GRF40_6_buffer[!clk]) ||(GRF40_7_buffer[clk] != GRF40_7_buffer[!clk]) ||(GRF40_8_buffer[clk] != GRF40_8_buffer[!clk]) ||(GRF40_9_buffer[clk] != GRF40_9_buffer[!clk]) ||(GRF40_10_buffer[clk] != GRF40_10_buffer[!clk]) ||(GRF40_11_buffer[clk] != GRF40_11_buffer[!clk]) ||(GRF40_12_buffer[clk] != GRF40_12_buffer[!clk]) ||(GRF40_13_buffer[clk] != GRF40_13_buffer[!clk]) ||(GRF40_14_buffer[clk] != GRF40_14_buffer[!clk]) ||(GRF40_15_buffer[clk] != GRF40_15_buffer[!clk]) ||(GRF40_16_buffer[clk] != GRF40_16_buffer[!clk]) ||(GRF40_17_buffer[clk] != GRF40_17_buffer[!clk]) ||(GRF40_18_buffer[clk] != GRF40_18_buffer[!clk]) ||(GRF40_19_buffer[clk] != GRF40_19_buffer[!clk]) ||(GRF40_20_buffer[clk] != GRF40_20_buffer[!clk]) ||(GRF40_21_buffer[clk] != GRF40_21_buffer[!clk]) ||(GRF40_22_buffer[clk] != GRF40_22_buffer[!clk]) ||(GRF40_23_buffer[clk] != GRF40_23_buffer[!clk]) ||(GRF40_24_buffer[clk] != GRF40_24_buffer[!clk]) ||(GRF40_25_buffer[clk] != GRF40_25_buffer[!clk]) ||(GRF40_26_buffer[clk] != GRF40_26_buffer[!clk]) ||(GRF40_27_buffer[clk] != GRF40_27_buffer[!clk]) ||(GRF40_28_buffer[clk] != GRF40_28_buffer[!clk]) ||(GRF40_29_buffer[clk] != GRF40_29_buffer[!clk]) ||(GRF40_30_buffer[clk] != GRF40_30_buffer[!clk]) ||(GRF40_31_buffer[clk] != GRF40_31_buffer[!clk]) ||(GRF48_0_buffer[clk] != GRF48_0_buffer[!clk]) ||(GRF48_1_buffer[clk] != GRF48_1_buffer[!clk]) ||(GRF48_2_buffer[clk] != GRF48_2_buffer[!clk]) ||(GRF48_3_buffer[clk] != GRF48_3_buffer[!clk]) ||(GRF48_4_buffer[clk] != GRF48_4_buffer[!clk]) ||(GRF48_5_buffer[clk] != GRF48_5_buffer[!clk]) ||(GRF48_6_buffer[clk] != GRF48_6_buffer[!clk]) ||(GRF48_7_buffer[clk] != GRF48_7_buffer[!clk]) ||(GRF48_8_buffer[clk] != GRF48_8_buffer[!clk]) ||(GRF48_9_buffer[clk] != GRF48_9_buffer[!clk]) ||(GRF48_10_buffer[clk] != GRF48_10_buffer[!clk]) ||(GRF48_11_buffer[clk] != GRF48_11_buffer[!clk]) ||(GRF48_12_buffer[clk] != GRF48_12_buffer[!clk]) ||(GRF48_13_buffer[clk] != GRF48_13_buffer[!clk]) ||(GRF48_14_buffer[clk] != GRF48_14_buffer[!clk]) ||(GRF48_15_buffer[clk] != GRF48_15_buffer[!clk]) ||(GRF48_16_buffer[clk] != GRF48_16_buffer[!clk]) ||(GRF48_17_buffer[clk] != GRF48_17_buffer[!clk]) ||(GRF48_18_buffer[clk] != GRF48_18_buffer[!clk]) ||(GRF48_19_buffer[clk] != GRF48_19_buffer[!clk]) ||(GRF48_20_buffer[clk] != GRF48_20_buffer[!clk]) ||(GRF48_21_buffer[clk] != GRF48_21_buffer[!clk]) ||(GRF48_22_buffer[clk] != GRF48_22_buffer[!clk]) ||(GRF48_23_buffer[clk] != GRF48_23_buffer[!clk]) ||(GRF48_24_buffer[clk] != GRF48_24_buffer[!clk]) ||(GRF48_25_buffer[clk] != GRF48_25_buffer[!clk]) ||(GRF48_26_buffer[clk] != GRF48_26_buffer[!clk]) ||(GRF48_27_buffer[clk] != GRF48_27_buffer[!clk]) ||(GRF48_28_buffer[clk] != GRF48_28_buffer[!clk]) ||(GRF48_29_buffer[clk] != GRF48_29_buffer[!clk]) ||(GRF48_30_buffer[clk] != GRF48_30_buffer[!clk]) ||(GRF48_31_buffer[clk] != GRF48_31_buffer[!clk]) ||(GRF56_0_buffer[clk] != GRF56_0_buffer[!clk]) ||(GRF56_1_buffer[clk] != GRF56_1_buffer[!clk]) ||(GRF56_2_buffer[clk] != GRF56_2_buffer[!clk]) ||(GRF56_3_buffer[clk] != GRF56_3_buffer[!clk]) ||(GRF56_4_buffer[clk] != GRF56_4_buffer[!clk]) ||(GRF56_5_buffer[clk] != GRF56_5_buffer[!clk]) ||(GRF56_6_buffer[clk] != GRF56_6_buffer[!clk]) ||(GRF56_7_buffer[clk] != GRF56_7_buffer[!clk]) ||(GRF56_8_buffer[clk] != GRF56_8_buffer[!clk]) ||(GRF56_9_buffer[clk] != GRF56_9_buffer[!clk]) ||(GRF56_10_buffer[clk] != GRF56_10_buffer[!clk]) ||(GRF56_11_buffer[clk] != GRF56_11_buffer[!clk]) ||(GRF56_12_buffer[clk] != GRF56_12_buffer[!clk]) ||(GRF56_13_buffer[clk] != GRF56_13_buffer[!clk]) ||(GRF56_14_buffer[clk] != GRF56_14_buffer[!clk]) ||(GRF56_15_buffer[clk] != GRF56_15_buffer[!clk]) ||(GRF56_16_buffer[clk] != GRF56_16_buffer[!clk]) ||(GRF56_17_buffer[clk] != GRF56_17_buffer[!clk]) ||(GRF56_18_buffer[clk] != GRF56_18_buffer[!clk]) ||(GRF56_19_buffer[clk] != GRF56_19_buffer[!clk]) ||(GRF56_20_buffer[clk] != GRF56_20_buffer[!clk]) ||(GRF56_21_buffer[clk] != GRF56_21_buffer[!clk]) ||(GRF56_22_buffer[clk] != GRF56_22_buffer[!clk]) ||(GRF56_23_buffer[clk] != GRF56_23_buffer[!clk]) ||(GRF56_24_buffer[clk] != GRF56_24_buffer[!clk]) ||(GRF56_25_buffer[clk] != GRF56_25_buffer[!clk]) ||(GRF56_26_buffer[clk] != GRF56_26_buffer[!clk]) ||(GRF56_27_buffer[clk] != GRF56_27_buffer[!clk]) ||(GRF56_28_buffer[clk] != GRF56_28_buffer[!clk]) ||(GRF56_29_buffer[clk] != GRF56_29_buffer[!clk]) ||(GRF56_30_buffer[clk] != GRF56_30_buffer[!clk]) ||(GRF56_31_buffer[clk] != GRF56_31_buffer[!clk]) ) begin
      warp0_sig = 1'b1;
    end else begin
      warp0_sig = 1'b0;
    end

    if ((GRF1_0_buffer[clk] != GRF1_0_buffer[!clk]) ||(GRF1_1_buffer[clk] != GRF1_1_buffer[!clk]) ||(GRF1_2_buffer[clk] != GRF1_2_buffer[!clk]) ||(GRF1_3_buffer[clk] != GRF1_3_buffer[!clk]) ||(GRF1_4_buffer[clk] != GRF1_4_buffer[!clk]) ||(GRF1_5_buffer[clk] != GRF1_5_buffer[!clk]) ||(GRF1_6_buffer[clk] != GRF1_6_buffer[!clk]) ||(GRF1_7_buffer[clk] != GRF1_7_buffer[!clk]) ||(GRF1_8_buffer[clk] != GRF1_8_buffer[!clk]) ||(GRF1_9_buffer[clk] != GRF1_9_buffer[!clk]) ||(GRF1_10_buffer[clk] != GRF1_10_buffer[!clk]) ||(GRF1_11_buffer[clk] != GRF1_11_buffer[!clk]) ||(GRF1_12_buffer[clk] != GRF1_12_buffer[!clk]) ||(GRF1_13_buffer[clk] != GRF1_13_buffer[!clk]) ||(GRF1_14_buffer[clk] != GRF1_14_buffer[!clk]) ||(GRF1_15_buffer[clk] != GRF1_15_buffer[!clk]) ||(GRF1_16_buffer[clk] != GRF1_16_buffer[!clk]) ||(GRF1_17_buffer[clk] != GRF1_17_buffer[!clk]) ||(GRF1_18_buffer[clk] != GRF1_18_buffer[!clk]) ||(GRF1_19_buffer[clk] != GRF1_19_buffer[!clk]) ||(GRF1_20_buffer[clk] != GRF1_20_buffer[!clk]) ||(GRF1_21_buffer[clk] != GRF1_21_buffer[!clk]) ||(GRF1_22_buffer[clk] != GRF1_22_buffer[!clk]) ||(GRF1_23_buffer[clk] != GRF1_23_buffer[!clk]) ||(GRF1_24_buffer[clk] != GRF1_24_buffer[!clk]) ||(GRF1_25_buffer[clk] != GRF1_25_buffer[!clk]) ||(GRF1_26_buffer[clk] != GRF1_26_buffer[!clk]) ||(GRF1_27_buffer[clk] != GRF1_27_buffer[!clk]) ||(GRF1_28_buffer[clk] != GRF1_28_buffer[!clk]) ||(GRF1_29_buffer[clk] != GRF1_29_buffer[!clk]) ||(GRF1_30_buffer[clk] != GRF1_30_buffer[!clk]) ||(GRF1_31_buffer[clk] != GRF1_31_buffer[!clk]) ||(GRF9_0_buffer[clk] != GRF9_0_buffer[!clk]) ||(GRF9_1_buffer[clk] != GRF9_1_buffer[!clk]) ||(GRF9_2_buffer[clk] != GRF9_2_buffer[!clk]) ||(GRF9_3_buffer[clk] != GRF9_3_buffer[!clk]) ||(GRF9_4_buffer[clk] != GRF9_4_buffer[!clk]) ||(GRF9_5_buffer[clk] != GRF9_5_buffer[!clk]) ||(GRF9_6_buffer[clk] != GRF9_6_buffer[!clk]) ||(GRF9_7_buffer[clk] != GRF9_7_buffer[!clk]) ||(GRF9_8_buffer[clk] != GRF9_8_buffer[!clk]) ||(GRF9_9_buffer[clk] != GRF9_9_buffer[!clk]) ||(GRF9_10_buffer[clk] != GRF9_10_buffer[!clk]) ||(GRF9_11_buffer[clk] != GRF9_11_buffer[!clk]) ||(GRF9_12_buffer[clk] != GRF9_12_buffer[!clk]) ||(GRF9_13_buffer[clk] != GRF9_13_buffer[!clk]) ||(GRF9_14_buffer[clk] != GRF9_14_buffer[!clk]) ||(GRF9_15_buffer[clk] != GRF9_15_buffer[!clk]) ||(GRF9_16_buffer[clk] != GRF9_16_buffer[!clk]) ||(GRF9_17_buffer[clk] != GRF9_17_buffer[!clk]) ||(GRF9_18_buffer[clk] != GRF9_18_buffer[!clk]) ||(GRF9_19_buffer[clk] != GRF9_19_buffer[!clk]) ||(GRF9_20_buffer[clk] != GRF9_20_buffer[!clk]) ||(GRF9_21_buffer[clk] != GRF9_21_buffer[!clk]) ||(GRF9_22_buffer[clk] != GRF9_22_buffer[!clk]) ||(GRF9_23_buffer[clk] != GRF9_23_buffer[!clk]) ||(GRF9_24_buffer[clk] != GRF9_24_buffer[!clk]) ||(GRF9_25_buffer[clk] != GRF9_25_buffer[!clk]) ||(GRF9_26_buffer[clk] != GRF9_26_buffer[!clk]) ||(GRF9_27_buffer[clk] != GRF9_27_buffer[!clk]) ||(GRF9_28_buffer[clk] != GRF9_28_buffer[!clk]) ||(GRF9_29_buffer[clk] != GRF9_29_buffer[!clk]) ||(GRF9_30_buffer[clk] != GRF9_30_buffer[!clk]) ||(GRF9_31_buffer[clk] != GRF9_31_buffer[!clk]) ||(GRF17_0_buffer[clk] != GRF17_0_buffer[!clk]) ||(GRF17_1_buffer[clk] != GRF17_1_buffer[!clk]) ||(GRF17_2_buffer[clk] != GRF17_2_buffer[!clk]) ||(GRF17_3_buffer[clk] != GRF17_3_buffer[!clk]) ||(GRF17_4_buffer[clk] != GRF17_4_buffer[!clk]) ||(GRF17_5_buffer[clk] != GRF17_5_buffer[!clk]) ||(GRF17_6_buffer[clk] != GRF17_6_buffer[!clk]) ||(GRF17_7_buffer[clk] != GRF17_7_buffer[!clk]) ||(GRF17_8_buffer[clk] != GRF17_8_buffer[!clk]) ||(GRF17_9_buffer[clk] != GRF17_9_buffer[!clk]) ||(GRF17_10_buffer[clk] != GRF17_10_buffer[!clk]) ||(GRF17_11_buffer[clk] != GRF17_11_buffer[!clk]) ||(GRF17_12_buffer[clk] != GRF17_12_buffer[!clk]) ||(GRF17_13_buffer[clk] != GRF17_13_buffer[!clk]) ||(GRF17_14_buffer[clk] != GRF17_14_buffer[!clk]) ||(GRF17_15_buffer[clk] != GRF17_15_buffer[!clk]) ||(GRF17_16_buffer[clk] != GRF17_16_buffer[!clk]) ||(GRF17_17_buffer[clk] != GRF17_17_buffer[!clk]) ||(GRF17_18_buffer[clk] != GRF17_18_buffer[!clk]) ||(GRF17_19_buffer[clk] != GRF17_19_buffer[!clk]) ||(GRF17_20_buffer[clk] != GRF17_20_buffer[!clk]) ||(GRF17_21_buffer[clk] != GRF17_21_buffer[!clk]) ||(GRF17_22_buffer[clk] != GRF17_22_buffer[!clk]) ||(GRF17_23_buffer[clk] != GRF17_23_buffer[!clk]) ||(GRF17_24_buffer[clk] != GRF17_24_buffer[!clk]) ||(GRF17_25_buffer[clk] != GRF17_25_buffer[!clk]) ||(GRF17_26_buffer[clk] != GRF17_26_buffer[!clk]) ||(GRF17_27_buffer[clk] != GRF17_27_buffer[!clk]) ||(GRF17_28_buffer[clk] != GRF17_28_buffer[!clk]) ||(GRF17_29_buffer[clk] != GRF17_29_buffer[!clk]) ||(GRF17_30_buffer[clk] != GRF17_30_buffer[!clk]) ||(GRF17_31_buffer[clk] != GRF17_31_buffer[!clk]) ||(GRF25_0_buffer[clk] != GRF25_0_buffer[!clk]) ||(GRF25_1_buffer[clk] != GRF25_1_buffer[!clk]) ||(GRF25_2_buffer[clk] != GRF25_2_buffer[!clk]) ||(GRF25_3_buffer[clk] != GRF25_3_buffer[!clk]) ||(GRF25_4_buffer[clk] != GRF25_4_buffer[!clk]) ||(GRF25_5_buffer[clk] != GRF25_5_buffer[!clk]) ||(GRF25_6_buffer[clk] != GRF25_6_buffer[!clk]) ||(GRF25_7_buffer[clk] != GRF25_7_buffer[!clk]) ||(GRF25_8_buffer[clk] != GRF25_8_buffer[!clk]) ||(GRF25_9_buffer[clk] != GRF25_9_buffer[!clk]) ||(GRF25_10_buffer[clk] != GRF25_10_buffer[!clk]) ||(GRF25_11_buffer[clk] != GRF25_11_buffer[!clk]) ||(GRF25_12_buffer[clk] != GRF25_12_buffer[!clk]) ||(GRF25_13_buffer[clk] != GRF25_13_buffer[!clk]) ||(GRF25_14_buffer[clk] != GRF25_14_buffer[!clk]) ||(GRF25_15_buffer[clk] != GRF25_15_buffer[!clk]) ||(GRF25_16_buffer[clk] != GRF25_16_buffer[!clk]) ||(GRF25_17_buffer[clk] != GRF25_17_buffer[!clk]) ||(GRF25_18_buffer[clk] != GRF25_18_buffer[!clk]) ||(GRF25_19_buffer[clk] != GRF25_19_buffer[!clk]) ||(GRF25_20_buffer[clk] != GRF25_20_buffer[!clk]) ||(GRF25_21_buffer[clk] != GRF25_21_buffer[!clk]) ||(GRF25_22_buffer[clk] != GRF25_22_buffer[!clk]) ||(GRF25_23_buffer[clk] != GRF25_23_buffer[!clk]) ||(GRF25_24_buffer[clk] != GRF25_24_buffer[!clk]) ||(GRF25_25_buffer[clk] != GRF25_25_buffer[!clk]) ||(GRF25_26_buffer[clk] != GRF25_26_buffer[!clk]) ||(GRF25_27_buffer[clk] != GRF25_27_buffer[!clk]) ||(GRF25_28_buffer[clk] != GRF25_28_buffer[!clk]) ||(GRF25_29_buffer[clk] != GRF25_29_buffer[!clk]) ||(GRF25_30_buffer[clk] != GRF25_30_buffer[!clk]) ||(GRF25_31_buffer[clk] != GRF25_31_buffer[!clk]) ||(GRF33_0_buffer[clk] != GRF33_0_buffer[!clk]) ||(GRF33_1_buffer[clk] != GRF33_1_buffer[!clk]) ||(GRF33_2_buffer[clk] != GRF33_2_buffer[!clk]) ||(GRF33_3_buffer[clk] != GRF33_3_buffer[!clk]) ||(GRF33_4_buffer[clk] != GRF33_4_buffer[!clk]) ||(GRF33_5_buffer[clk] != GRF33_5_buffer[!clk]) ||(GRF33_6_buffer[clk] != GRF33_6_buffer[!clk]) ||(GRF33_7_buffer[clk] != GRF33_7_buffer[!clk]) ||(GRF33_8_buffer[clk] != GRF33_8_buffer[!clk]) ||(GRF33_9_buffer[clk] != GRF33_9_buffer[!clk]) ||(GRF33_10_buffer[clk] != GRF33_10_buffer[!clk]) ||(GRF33_11_buffer[clk] != GRF33_11_buffer[!clk]) ||(GRF33_12_buffer[clk] != GRF33_12_buffer[!clk]) ||(GRF33_13_buffer[clk] != GRF33_13_buffer[!clk]) ||(GRF33_14_buffer[clk] != GRF33_14_buffer[!clk]) ||(GRF33_15_buffer[clk] != GRF33_15_buffer[!clk]) ||(GRF33_16_buffer[clk] != GRF33_16_buffer[!clk]) ||(GRF33_17_buffer[clk] != GRF33_17_buffer[!clk]) ||(GRF33_18_buffer[clk] != GRF33_18_buffer[!clk]) ||(GRF33_19_buffer[clk] != GRF33_19_buffer[!clk]) ||(GRF33_20_buffer[clk] != GRF33_20_buffer[!clk]) ||(GRF33_21_buffer[clk] != GRF33_21_buffer[!clk]) ||(GRF33_22_buffer[clk] != GRF33_22_buffer[!clk]) ||(GRF33_23_buffer[clk] != GRF33_23_buffer[!clk]) ||(GRF33_24_buffer[clk] != GRF33_24_buffer[!clk]) ||(GRF33_25_buffer[clk] != GRF33_25_buffer[!clk]) ||(GRF33_26_buffer[clk] != GRF33_26_buffer[!clk]) ||(GRF33_27_buffer[clk] != GRF33_27_buffer[!clk]) ||(GRF33_28_buffer[clk] != GRF33_28_buffer[!clk]) ||(GRF33_29_buffer[clk] != GRF33_29_buffer[!clk]) ||(GRF33_30_buffer[clk] != GRF33_30_buffer[!clk]) ||(GRF33_31_buffer[clk] != GRF33_31_buffer[!clk]) ||(GRF41_0_buffer[clk] != GRF41_0_buffer[!clk]) ||(GRF41_1_buffer[clk] != GRF41_1_buffer[!clk]) ||(GRF41_2_buffer[clk] != GRF41_2_buffer[!clk]) ||(GRF41_3_buffer[clk] != GRF41_3_buffer[!clk]) ||(GRF41_4_buffer[clk] != GRF41_4_buffer[!clk]) ||(GRF41_5_buffer[clk] != GRF41_5_buffer[!clk]) ||(GRF41_6_buffer[clk] != GRF41_6_buffer[!clk]) ||(GRF41_7_buffer[clk] != GRF41_7_buffer[!clk]) ||(GRF41_8_buffer[clk] != GRF41_8_buffer[!clk]) ||(GRF41_9_buffer[clk] != GRF41_9_buffer[!clk]) ||(GRF41_10_buffer[clk] != GRF41_10_buffer[!clk]) ||(GRF41_11_buffer[clk] != GRF41_11_buffer[!clk]) ||(GRF41_12_buffer[clk] != GRF41_12_buffer[!clk]) ||(GRF41_13_buffer[clk] != GRF41_13_buffer[!clk]) ||(GRF41_14_buffer[clk] != GRF41_14_buffer[!clk]) ||(GRF41_15_buffer[clk] != GRF41_15_buffer[!clk]) ||(GRF41_16_buffer[clk] != GRF41_16_buffer[!clk]) ||(GRF41_17_buffer[clk] != GRF41_17_buffer[!clk]) ||(GRF41_18_buffer[clk] != GRF41_18_buffer[!clk]) ||(GRF41_19_buffer[clk] != GRF41_19_buffer[!clk]) ||(GRF41_20_buffer[clk] != GRF41_20_buffer[!clk]) ||(GRF41_21_buffer[clk] != GRF41_21_buffer[!clk]) ||(GRF41_22_buffer[clk] != GRF41_22_buffer[!clk]) ||(GRF41_23_buffer[clk] != GRF41_23_buffer[!clk]) ||(GRF41_24_buffer[clk] != GRF41_24_buffer[!clk]) ||(GRF41_25_buffer[clk] != GRF41_25_buffer[!clk]) ||(GRF41_26_buffer[clk] != GRF41_26_buffer[!clk]) ||(GRF41_27_buffer[clk] != GRF41_27_buffer[!clk]) ||(GRF41_28_buffer[clk] != GRF41_28_buffer[!clk]) ||(GRF41_29_buffer[clk] != GRF41_29_buffer[!clk]) ||(GRF41_30_buffer[clk] != GRF41_30_buffer[!clk]) ||(GRF41_31_buffer[clk] != GRF41_31_buffer[!clk]) ||(GRF49_0_buffer[clk] != GRF49_0_buffer[!clk]) ||(GRF49_1_buffer[clk] != GRF49_1_buffer[!clk]) ||(GRF49_2_buffer[clk] != GRF49_2_buffer[!clk]) ||(GRF49_3_buffer[clk] != GRF49_3_buffer[!clk]) ||(GRF49_4_buffer[clk] != GRF49_4_buffer[!clk]) ||(GRF49_5_buffer[clk] != GRF49_5_buffer[!clk]) ||(GRF49_6_buffer[clk] != GRF49_6_buffer[!clk]) ||(GRF49_7_buffer[clk] != GRF49_7_buffer[!clk]) ||(GRF49_8_buffer[clk] != GRF49_8_buffer[!clk]) ||(GRF49_9_buffer[clk] != GRF49_9_buffer[!clk]) ||(GRF49_10_buffer[clk] != GRF49_10_buffer[!clk]) ||(GRF49_11_buffer[clk] != GRF49_11_buffer[!clk]) ||(GRF49_12_buffer[clk] != GRF49_12_buffer[!clk]) ||(GRF49_13_buffer[clk] != GRF49_13_buffer[!clk]) ||(GRF49_14_buffer[clk] != GRF49_14_buffer[!clk]) ||(GRF49_15_buffer[clk] != GRF49_15_buffer[!clk]) ||(GRF49_16_buffer[clk] != GRF49_16_buffer[!clk]) ||(GRF49_17_buffer[clk] != GRF49_17_buffer[!clk]) ||(GRF49_18_buffer[clk] != GRF49_18_buffer[!clk]) ||(GRF49_19_buffer[clk] != GRF49_19_buffer[!clk]) ||(GRF49_20_buffer[clk] != GRF49_20_buffer[!clk]) ||(GRF49_21_buffer[clk] != GRF49_21_buffer[!clk]) ||(GRF49_22_buffer[clk] != GRF49_22_buffer[!clk]) ||(GRF49_23_buffer[clk] != GRF49_23_buffer[!clk]) ||(GRF49_24_buffer[clk] != GRF49_24_buffer[!clk]) ||(GRF49_25_buffer[clk] != GRF49_25_buffer[!clk]) ||(GRF49_26_buffer[clk] != GRF49_26_buffer[!clk]) ||(GRF49_27_buffer[clk] != GRF49_27_buffer[!clk]) ||(GRF49_28_buffer[clk] != GRF49_28_buffer[!clk]) ||(GRF49_29_buffer[clk] != GRF49_29_buffer[!clk]) ||(GRF49_30_buffer[clk] != GRF49_30_buffer[!clk]) ||(GRF49_31_buffer[clk] != GRF49_31_buffer[!clk]) ||(GRF57_0_buffer[clk] != GRF57_0_buffer[!clk]) ||(GRF57_1_buffer[clk] != GRF57_1_buffer[!clk]) ||(GRF57_2_buffer[clk] != GRF57_2_buffer[!clk]) ||(GRF57_3_buffer[clk] != GRF57_3_buffer[!clk]) ||(GRF57_4_buffer[clk] != GRF57_4_buffer[!clk]) ||(GRF57_5_buffer[clk] != GRF57_5_buffer[!clk]) ||(GRF57_6_buffer[clk] != GRF57_6_buffer[!clk]) ||(GRF57_7_buffer[clk] != GRF57_7_buffer[!clk]) ||(GRF57_8_buffer[clk] != GRF57_8_buffer[!clk]) ||(GRF57_9_buffer[clk] != GRF57_9_buffer[!clk]) ||(GRF57_10_buffer[clk] != GRF57_10_buffer[!clk]) ||(GRF57_11_buffer[clk] != GRF57_11_buffer[!clk]) ||(GRF57_12_buffer[clk] != GRF57_12_buffer[!clk]) ||(GRF57_13_buffer[clk] != GRF57_13_buffer[!clk]) ||(GRF57_14_buffer[clk] != GRF57_14_buffer[!clk]) ||(GRF57_15_buffer[clk] != GRF57_15_buffer[!clk]) ||(GRF57_16_buffer[clk] != GRF57_16_buffer[!clk]) ||(GRF57_17_buffer[clk] != GRF57_17_buffer[!clk]) ||(GRF57_18_buffer[clk] != GRF57_18_buffer[!clk]) ||(GRF57_19_buffer[clk] != GRF57_19_buffer[!clk]) ||(GRF57_20_buffer[clk] != GRF57_20_buffer[!clk]) ||(GRF57_21_buffer[clk] != GRF57_21_buffer[!clk]) ||(GRF57_22_buffer[clk] != GRF57_22_buffer[!clk]) ||(GRF57_23_buffer[clk] != GRF57_23_buffer[!clk]) ||(GRF57_24_buffer[clk] != GRF57_24_buffer[!clk]) ||(GRF57_25_buffer[clk] != GRF57_25_buffer[!clk]) ||(GRF57_26_buffer[clk] != GRF57_26_buffer[!clk]) ||(GRF57_27_buffer[clk] != GRF57_27_buffer[!clk]) ||(GRF57_28_buffer[clk] != GRF57_28_buffer[!clk]) ||(GRF57_29_buffer[clk] != GRF57_29_buffer[!clk]) ||(GRF57_30_buffer[clk] != GRF57_30_buffer[!clk]) ||(GRF57_31_buffer[clk] != GRF57_31_buffer[!clk]) ) begin
      warp1_sig = 1'b1;
    end else begin
      warp1_sig = 1'b0;
    end

    if ((GRF2_0_buffer[clk] != GRF2_0_buffer[!clk]) ||(GRF2_1_buffer[clk] != GRF2_1_buffer[!clk]) ||(GRF2_2_buffer[clk] != GRF2_2_buffer[!clk]) ||(GRF2_3_buffer[clk] != GRF2_3_buffer[!clk]) ||(GRF2_4_buffer[clk] != GRF2_4_buffer[!clk]) ||(GRF2_5_buffer[clk] != GRF2_5_buffer[!clk]) ||(GRF2_6_buffer[clk] != GRF2_6_buffer[!clk]) ||(GRF2_7_buffer[clk] != GRF2_7_buffer[!clk]) ||(GRF2_8_buffer[clk] != GRF2_8_buffer[!clk]) ||(GRF2_9_buffer[clk] != GRF2_9_buffer[!clk]) ||(GRF2_10_buffer[clk] != GRF2_10_buffer[!clk]) ||(GRF2_11_buffer[clk] != GRF2_11_buffer[!clk]) ||(GRF2_12_buffer[clk] != GRF2_12_buffer[!clk]) ||(GRF2_13_buffer[clk] != GRF2_13_buffer[!clk]) ||(GRF2_14_buffer[clk] != GRF2_14_buffer[!clk]) ||(GRF2_15_buffer[clk] != GRF2_15_buffer[!clk]) ||(GRF2_16_buffer[clk] != GRF2_16_buffer[!clk]) ||(GRF2_17_buffer[clk] != GRF2_17_buffer[!clk]) ||(GRF2_18_buffer[clk] != GRF2_18_buffer[!clk]) ||(GRF2_19_buffer[clk] != GRF2_19_buffer[!clk]) ||(GRF2_20_buffer[clk] != GRF2_20_buffer[!clk]) ||(GRF2_21_buffer[clk] != GRF2_21_buffer[!clk]) ||(GRF2_22_buffer[clk] != GRF2_22_buffer[!clk]) ||(GRF2_23_buffer[clk] != GRF2_23_buffer[!clk]) ||(GRF2_24_buffer[clk] != GRF2_24_buffer[!clk]) ||(GRF2_25_buffer[clk] != GRF2_25_buffer[!clk]) ||(GRF2_26_buffer[clk] != GRF2_26_buffer[!clk]) ||(GRF2_27_buffer[clk] != GRF2_27_buffer[!clk]) ||(GRF2_28_buffer[clk] != GRF2_28_buffer[!clk]) ||(GRF2_29_buffer[clk] != GRF2_29_buffer[!clk]) ||(GRF2_30_buffer[clk] != GRF2_30_buffer[!clk]) ||(GRF2_31_buffer[clk] != GRF2_31_buffer[!clk]) ||(GRF10_0_buffer[clk] != GRF10_0_buffer[!clk]) ||(GRF10_1_buffer[clk] != GRF10_1_buffer[!clk]) ||(GRF10_2_buffer[clk] != GRF10_2_buffer[!clk]) ||(GRF10_3_buffer[clk] != GRF10_3_buffer[!clk]) ||(GRF10_4_buffer[clk] != GRF10_4_buffer[!clk]) ||(GRF10_5_buffer[clk] != GRF10_5_buffer[!clk]) ||(GRF10_6_buffer[clk] != GRF10_6_buffer[!clk]) ||(GRF10_7_buffer[clk] != GRF10_7_buffer[!clk]) ||(GRF10_8_buffer[clk] != GRF10_8_buffer[!clk]) ||(GRF10_9_buffer[clk] != GRF10_9_buffer[!clk]) ||(GRF10_10_buffer[clk] != GRF10_10_buffer[!clk]) ||(GRF10_11_buffer[clk] != GRF10_11_buffer[!clk]) ||(GRF10_12_buffer[clk] != GRF10_12_buffer[!clk]) ||(GRF10_13_buffer[clk] != GRF10_13_buffer[!clk]) ||(GRF10_14_buffer[clk] != GRF10_14_buffer[!clk]) ||(GRF10_15_buffer[clk] != GRF10_15_buffer[!clk]) ||(GRF10_16_buffer[clk] != GRF10_16_buffer[!clk]) ||(GRF10_17_buffer[clk] != GRF10_17_buffer[!clk]) ||(GRF10_18_buffer[clk] != GRF10_18_buffer[!clk]) ||(GRF10_19_buffer[clk] != GRF10_19_buffer[!clk]) ||(GRF10_20_buffer[clk] != GRF10_20_buffer[!clk]) ||(GRF10_21_buffer[clk] != GRF10_21_buffer[!clk]) ||(GRF10_22_buffer[clk] != GRF10_22_buffer[!clk]) ||(GRF10_23_buffer[clk] != GRF10_23_buffer[!clk]) ||(GRF10_24_buffer[clk] != GRF10_24_buffer[!clk]) ||(GRF10_25_buffer[clk] != GRF10_25_buffer[!clk]) ||(GRF10_26_buffer[clk] != GRF10_26_buffer[!clk]) ||(GRF10_27_buffer[clk] != GRF10_27_buffer[!clk]) ||(GRF10_28_buffer[clk] != GRF10_28_buffer[!clk]) ||(GRF10_29_buffer[clk] != GRF10_29_buffer[!clk]) ||(GRF10_30_buffer[clk] != GRF10_30_buffer[!clk]) ||(GRF10_31_buffer[clk] != GRF10_31_buffer[!clk]) ||(GRF18_0_buffer[clk] != GRF18_0_buffer[!clk]) ||(GRF18_1_buffer[clk] != GRF18_1_buffer[!clk]) ||(GRF18_2_buffer[clk] != GRF18_2_buffer[!clk]) ||(GRF18_3_buffer[clk] != GRF18_3_buffer[!clk]) ||(GRF18_4_buffer[clk] != GRF18_4_buffer[!clk]) ||(GRF18_5_buffer[clk] != GRF18_5_buffer[!clk]) ||(GRF18_6_buffer[clk] != GRF18_6_buffer[!clk]) ||(GRF18_7_buffer[clk] != GRF18_7_buffer[!clk]) ||(GRF18_8_buffer[clk] != GRF18_8_buffer[!clk]) ||(GRF18_9_buffer[clk] != GRF18_9_buffer[!clk]) ||(GRF18_10_buffer[clk] != GRF18_10_buffer[!clk]) ||(GRF18_11_buffer[clk] != GRF18_11_buffer[!clk]) ||(GRF18_12_buffer[clk] != GRF18_12_buffer[!clk]) ||(GRF18_13_buffer[clk] != GRF18_13_buffer[!clk]) ||(GRF18_14_buffer[clk] != GRF18_14_buffer[!clk]) ||(GRF18_15_buffer[clk] != GRF18_15_buffer[!clk]) ||(GRF18_16_buffer[clk] != GRF18_16_buffer[!clk]) ||(GRF18_17_buffer[clk] != GRF18_17_buffer[!clk]) ||(GRF18_18_buffer[clk] != GRF18_18_buffer[!clk]) ||(GRF18_19_buffer[clk] != GRF18_19_buffer[!clk]) ||(GRF18_20_buffer[clk] != GRF18_20_buffer[!clk]) ||(GRF18_21_buffer[clk] != GRF18_21_buffer[!clk]) ||(GRF18_22_buffer[clk] != GRF18_22_buffer[!clk]) ||(GRF18_23_buffer[clk] != GRF18_23_buffer[!clk]) ||(GRF18_24_buffer[clk] != GRF18_24_buffer[!clk]) ||(GRF18_25_buffer[clk] != GRF18_25_buffer[!clk]) ||(GRF18_26_buffer[clk] != GRF18_26_buffer[!clk]) ||(GRF18_27_buffer[clk] != GRF18_27_buffer[!clk]) ||(GRF18_28_buffer[clk] != GRF18_28_buffer[!clk]) ||(GRF18_29_buffer[clk] != GRF18_29_buffer[!clk]) ||(GRF18_30_buffer[clk] != GRF18_30_buffer[!clk]) ||(GRF18_31_buffer[clk] != GRF18_31_buffer[!clk]) ||(GRF26_0_buffer[clk] != GRF26_0_buffer[!clk]) ||(GRF26_1_buffer[clk] != GRF26_1_buffer[!clk]) ||(GRF26_2_buffer[clk] != GRF26_2_buffer[!clk]) ||(GRF26_3_buffer[clk] != GRF26_3_buffer[!clk]) ||(GRF26_4_buffer[clk] != GRF26_4_buffer[!clk]) ||(GRF26_5_buffer[clk] != GRF26_5_buffer[!clk]) ||(GRF26_6_buffer[clk] != GRF26_6_buffer[!clk]) ||(GRF26_7_buffer[clk] != GRF26_7_buffer[!clk]) ||(GRF26_8_buffer[clk] != GRF26_8_buffer[!clk]) ||(GRF26_9_buffer[clk] != GRF26_9_buffer[!clk]) ||(GRF26_10_buffer[clk] != GRF26_10_buffer[!clk]) ||(GRF26_11_buffer[clk] != GRF26_11_buffer[!clk]) ||(GRF26_12_buffer[clk] != GRF26_12_buffer[!clk]) ||(GRF26_13_buffer[clk] != GRF26_13_buffer[!clk]) ||(GRF26_14_buffer[clk] != GRF26_14_buffer[!clk]) ||(GRF26_15_buffer[clk] != GRF26_15_buffer[!clk]) ||(GRF26_16_buffer[clk] != GRF26_16_buffer[!clk]) ||(GRF26_17_buffer[clk] != GRF26_17_buffer[!clk]) ||(GRF26_18_buffer[clk] != GRF26_18_buffer[!clk]) ||(GRF26_19_buffer[clk] != GRF26_19_buffer[!clk]) ||(GRF26_20_buffer[clk] != GRF26_20_buffer[!clk]) ||(GRF26_21_buffer[clk] != GRF26_21_buffer[!clk]) ||(GRF26_22_buffer[clk] != GRF26_22_buffer[!clk]) ||(GRF26_23_buffer[clk] != GRF26_23_buffer[!clk]) ||(GRF26_24_buffer[clk] != GRF26_24_buffer[!clk]) ||(GRF26_25_buffer[clk] != GRF26_25_buffer[!clk]) ||(GRF26_26_buffer[clk] != GRF26_26_buffer[!clk]) ||(GRF26_27_buffer[clk] != GRF26_27_buffer[!clk]) ||(GRF26_28_buffer[clk] != GRF26_28_buffer[!clk]) ||(GRF26_29_buffer[clk] != GRF26_29_buffer[!clk]) ||(GRF26_30_buffer[clk] != GRF26_30_buffer[!clk]) ||(GRF26_31_buffer[clk] != GRF26_31_buffer[!clk]) ||(GRF34_0_buffer[clk] != GRF34_0_buffer[!clk]) ||(GRF34_1_buffer[clk] != GRF34_1_buffer[!clk]) ||(GRF34_2_buffer[clk] != GRF34_2_buffer[!clk]) ||(GRF34_3_buffer[clk] != GRF34_3_buffer[!clk]) ||(GRF34_4_buffer[clk] != GRF34_4_buffer[!clk]) ||(GRF34_5_buffer[clk] != GRF34_5_buffer[!clk]) ||(GRF34_6_buffer[clk] != GRF34_6_buffer[!clk]) ||(GRF34_7_buffer[clk] != GRF34_7_buffer[!clk]) ||(GRF34_8_buffer[clk] != GRF34_8_buffer[!clk]) ||(GRF34_9_buffer[clk] != GRF34_9_buffer[!clk]) ||(GRF34_10_buffer[clk] != GRF34_10_buffer[!clk]) ||(GRF34_11_buffer[clk] != GRF34_11_buffer[!clk]) ||(GRF34_12_buffer[clk] != GRF34_12_buffer[!clk]) ||(GRF34_13_buffer[clk] != GRF34_13_buffer[!clk]) ||(GRF34_14_buffer[clk] != GRF34_14_buffer[!clk]) ||(GRF34_15_buffer[clk] != GRF34_15_buffer[!clk]) ||(GRF34_16_buffer[clk] != GRF34_16_buffer[!clk]) ||(GRF34_17_buffer[clk] != GRF34_17_buffer[!clk]) ||(GRF34_18_buffer[clk] != GRF34_18_buffer[!clk]) ||(GRF34_19_buffer[clk] != GRF34_19_buffer[!clk]) ||(GRF34_20_buffer[clk] != GRF34_20_buffer[!clk]) ||(GRF34_21_buffer[clk] != GRF34_21_buffer[!clk]) ||(GRF34_22_buffer[clk] != GRF34_22_buffer[!clk]) ||(GRF34_23_buffer[clk] != GRF34_23_buffer[!clk]) ||(GRF34_24_buffer[clk] != GRF34_24_buffer[!clk]) ||(GRF34_25_buffer[clk] != GRF34_25_buffer[!clk]) ||(GRF34_26_buffer[clk] != GRF34_26_buffer[!clk]) ||(GRF34_27_buffer[clk] != GRF34_27_buffer[!clk]) ||(GRF34_28_buffer[clk] != GRF34_28_buffer[!clk]) ||(GRF34_29_buffer[clk] != GRF34_29_buffer[!clk]) ||(GRF34_30_buffer[clk] != GRF34_30_buffer[!clk]) ||(GRF34_31_buffer[clk] != GRF34_31_buffer[!clk]) ||(GRF42_0_buffer[clk] != GRF42_0_buffer[!clk]) ||(GRF42_1_buffer[clk] != GRF42_1_buffer[!clk]) ||(GRF42_2_buffer[clk] != GRF42_2_buffer[!clk]) ||(GRF42_3_buffer[clk] != GRF42_3_buffer[!clk]) ||(GRF42_4_buffer[clk] != GRF42_4_buffer[!clk]) ||(GRF42_5_buffer[clk] != GRF42_5_buffer[!clk]) ||(GRF42_6_buffer[clk] != GRF42_6_buffer[!clk]) ||(GRF42_7_buffer[clk] != GRF42_7_buffer[!clk]) ||(GRF42_8_buffer[clk] != GRF42_8_buffer[!clk]) ||(GRF42_9_buffer[clk] != GRF42_9_buffer[!clk]) ||(GRF42_10_buffer[clk] != GRF42_10_buffer[!clk]) ||(GRF42_11_buffer[clk] != GRF42_11_buffer[!clk]) ||(GRF42_12_buffer[clk] != GRF42_12_buffer[!clk]) ||(GRF42_13_buffer[clk] != GRF42_13_buffer[!clk]) ||(GRF42_14_buffer[clk] != GRF42_14_buffer[!clk]) ||(GRF42_15_buffer[clk] != GRF42_15_buffer[!clk]) ||(GRF42_16_buffer[clk] != GRF42_16_buffer[!clk]) ||(GRF42_17_buffer[clk] != GRF42_17_buffer[!clk]) ||(GRF42_18_buffer[clk] != GRF42_18_buffer[!clk]) ||(GRF42_19_buffer[clk] != GRF42_19_buffer[!clk]) ||(GRF42_20_buffer[clk] != GRF42_20_buffer[!clk]) ||(GRF42_21_buffer[clk] != GRF42_21_buffer[!clk]) ||(GRF42_22_buffer[clk] != GRF42_22_buffer[!clk]) ||(GRF42_23_buffer[clk] != GRF42_23_buffer[!clk]) ||(GRF42_24_buffer[clk] != GRF42_24_buffer[!clk]) ||(GRF42_25_buffer[clk] != GRF42_25_buffer[!clk]) ||(GRF42_26_buffer[clk] != GRF42_26_buffer[!clk]) ||(GRF42_27_buffer[clk] != GRF42_27_buffer[!clk]) ||(GRF42_28_buffer[clk] != GRF42_28_buffer[!clk]) ||(GRF42_29_buffer[clk] != GRF42_29_buffer[!clk]) ||(GRF42_30_buffer[clk] != GRF42_30_buffer[!clk]) ||(GRF42_31_buffer[clk] != GRF42_31_buffer[!clk]) ||(GRF50_0_buffer[clk] != GRF50_0_buffer[!clk]) ||(GRF50_1_buffer[clk] != GRF50_1_buffer[!clk]) ||(GRF50_2_buffer[clk] != GRF50_2_buffer[!clk]) ||(GRF50_3_buffer[clk] != GRF50_3_buffer[!clk]) ||(GRF50_4_buffer[clk] != GRF50_4_buffer[!clk]) ||(GRF50_5_buffer[clk] != GRF50_5_buffer[!clk]) ||(GRF50_6_buffer[clk] != GRF50_6_buffer[!clk]) ||(GRF50_7_buffer[clk] != GRF50_7_buffer[!clk]) ||(GRF50_8_buffer[clk] != GRF50_8_buffer[!clk]) ||(GRF50_9_buffer[clk] != GRF50_9_buffer[!clk]) ||(GRF50_10_buffer[clk] != GRF50_10_buffer[!clk]) ||(GRF50_11_buffer[clk] != GRF50_11_buffer[!clk]) ||(GRF50_12_buffer[clk] != GRF50_12_buffer[!clk]) ||(GRF50_13_buffer[clk] != GRF50_13_buffer[!clk]) ||(GRF50_14_buffer[clk] != GRF50_14_buffer[!clk]) ||(GRF50_15_buffer[clk] != GRF50_15_buffer[!clk]) ||(GRF50_16_buffer[clk] != GRF50_16_buffer[!clk]) ||(GRF50_17_buffer[clk] != GRF50_17_buffer[!clk]) ||(GRF50_18_buffer[clk] != GRF50_18_buffer[!clk]) ||(GRF50_19_buffer[clk] != GRF50_19_buffer[!clk]) ||(GRF50_20_buffer[clk] != GRF50_20_buffer[!clk]) ||(GRF50_21_buffer[clk] != GRF50_21_buffer[!clk]) ||(GRF50_22_buffer[clk] != GRF50_22_buffer[!clk]) ||(GRF50_23_buffer[clk] != GRF50_23_buffer[!clk]) ||(GRF50_24_buffer[clk] != GRF50_24_buffer[!clk]) ||(GRF50_25_buffer[clk] != GRF50_25_buffer[!clk]) ||(GRF50_26_buffer[clk] != GRF50_26_buffer[!clk]) ||(GRF50_27_buffer[clk] != GRF50_27_buffer[!clk]) ||(GRF50_28_buffer[clk] != GRF50_28_buffer[!clk]) ||(GRF50_29_buffer[clk] != GRF50_29_buffer[!clk]) ||(GRF50_30_buffer[clk] != GRF50_30_buffer[!clk]) ||(GRF50_31_buffer[clk] != GRF50_31_buffer[!clk]) ||(GRF58_0_buffer[clk] != GRF58_0_buffer[!clk]) ||(GRF58_1_buffer[clk] != GRF58_1_buffer[!clk]) ||(GRF58_2_buffer[clk] != GRF58_2_buffer[!clk]) ||(GRF58_3_buffer[clk] != GRF58_3_buffer[!clk]) ||(GRF58_4_buffer[clk] != GRF58_4_buffer[!clk]) ||(GRF58_5_buffer[clk] != GRF58_5_buffer[!clk]) ||(GRF58_6_buffer[clk] != GRF58_6_buffer[!clk]) ||(GRF58_7_buffer[clk] != GRF58_7_buffer[!clk]) ||(GRF58_8_buffer[clk] != GRF58_8_buffer[!clk]) ||(GRF58_9_buffer[clk] != GRF58_9_buffer[!clk]) ||(GRF58_10_buffer[clk] != GRF58_10_buffer[!clk]) ||(GRF58_11_buffer[clk] != GRF58_11_buffer[!clk]) ||(GRF58_12_buffer[clk] != GRF58_12_buffer[!clk]) ||(GRF58_13_buffer[clk] != GRF58_13_buffer[!clk]) ||(GRF58_14_buffer[clk] != GRF58_14_buffer[!clk]) ||(GRF58_15_buffer[clk] != GRF58_15_buffer[!clk]) ||(GRF58_16_buffer[clk] != GRF58_16_buffer[!clk]) ||(GRF58_17_buffer[clk] != GRF58_17_buffer[!clk]) ||(GRF58_18_buffer[clk] != GRF58_18_buffer[!clk]) ||(GRF58_19_buffer[clk] != GRF58_19_buffer[!clk]) ||(GRF58_20_buffer[clk] != GRF58_20_buffer[!clk]) ||(GRF58_21_buffer[clk] != GRF58_21_buffer[!clk]) ||(GRF58_22_buffer[clk] != GRF58_22_buffer[!clk]) ||(GRF58_23_buffer[clk] != GRF58_23_buffer[!clk]) ||(GRF58_24_buffer[clk] != GRF58_24_buffer[!clk]) ||(GRF58_25_buffer[clk] != GRF58_25_buffer[!clk]) ||(GRF58_26_buffer[clk] != GRF58_26_buffer[!clk]) ||(GRF58_27_buffer[clk] != GRF58_27_buffer[!clk]) ||(GRF58_28_buffer[clk] != GRF58_28_buffer[!clk]) ||(GRF58_29_buffer[clk] != GRF58_29_buffer[!clk]) ||(GRF58_30_buffer[clk] != GRF58_30_buffer[!clk]) ||(GRF58_31_buffer[clk] != GRF58_31_buffer[!clk]) ) begin
      warp2_sig = 1'b1;
    end else begin
      warp2_sig = 1'b0;
    end

    if ((GRF3_0_buffer[clk] != GRF3_0_buffer[!clk]) ||(GRF3_1_buffer[clk] != GRF3_1_buffer[!clk]) ||(GRF3_2_buffer[clk] != GRF3_2_buffer[!clk]) ||(GRF3_3_buffer[clk] != GRF3_3_buffer[!clk]) ||(GRF3_4_buffer[clk] != GRF3_4_buffer[!clk]) ||(GRF3_5_buffer[clk] != GRF3_5_buffer[!clk]) ||(GRF3_6_buffer[clk] != GRF3_6_buffer[!clk]) ||(GRF3_7_buffer[clk] != GRF3_7_buffer[!clk]) ||(GRF3_8_buffer[clk] != GRF3_8_buffer[!clk]) ||(GRF3_9_buffer[clk] != GRF3_9_buffer[!clk]) ||(GRF3_10_buffer[clk] != GRF3_10_buffer[!clk]) ||(GRF3_11_buffer[clk] != GRF3_11_buffer[!clk]) ||(GRF3_12_buffer[clk] != GRF3_12_buffer[!clk]) ||(GRF3_13_buffer[clk] != GRF3_13_buffer[!clk]) ||(GRF3_14_buffer[clk] != GRF3_14_buffer[!clk]) ||(GRF3_15_buffer[clk] != GRF3_15_buffer[!clk]) ||(GRF3_16_buffer[clk] != GRF3_16_buffer[!clk]) ||(GRF3_17_buffer[clk] != GRF3_17_buffer[!clk]) ||(GRF3_18_buffer[clk] != GRF3_18_buffer[!clk]) ||(GRF3_19_buffer[clk] != GRF3_19_buffer[!clk]) ||(GRF3_20_buffer[clk] != GRF3_20_buffer[!clk]) ||(GRF3_21_buffer[clk] != GRF3_21_buffer[!clk]) ||(GRF3_22_buffer[clk] != GRF3_22_buffer[!clk]) ||(GRF3_23_buffer[clk] != GRF3_23_buffer[!clk]) ||(GRF3_24_buffer[clk] != GRF3_24_buffer[!clk]) ||(GRF3_25_buffer[clk] != GRF3_25_buffer[!clk]) ||(GRF3_26_buffer[clk] != GRF3_26_buffer[!clk]) ||(GRF3_27_buffer[clk] != GRF3_27_buffer[!clk]) ||(GRF3_28_buffer[clk] != GRF3_28_buffer[!clk]) ||(GRF3_29_buffer[clk] != GRF3_29_buffer[!clk]) ||(GRF3_30_buffer[clk] != GRF3_30_buffer[!clk]) ||(GRF3_31_buffer[clk] != GRF3_31_buffer[!clk]) ||(GRF11_0_buffer[clk] != GRF11_0_buffer[!clk]) ||(GRF11_1_buffer[clk] != GRF11_1_buffer[!clk]) ||(GRF11_2_buffer[clk] != GRF11_2_buffer[!clk]) ||(GRF11_3_buffer[clk] != GRF11_3_buffer[!clk]) ||(GRF11_4_buffer[clk] != GRF11_4_buffer[!clk]) ||(GRF11_5_buffer[clk] != GRF11_5_buffer[!clk]) ||(GRF11_6_buffer[clk] != GRF11_6_buffer[!clk]) ||(GRF11_7_buffer[clk] != GRF11_7_buffer[!clk]) ||(GRF11_8_buffer[clk] != GRF11_8_buffer[!clk]) ||(GRF11_9_buffer[clk] != GRF11_9_buffer[!clk]) ||(GRF11_10_buffer[clk] != GRF11_10_buffer[!clk]) ||(GRF11_11_buffer[clk] != GRF11_11_buffer[!clk]) ||(GRF11_12_buffer[clk] != GRF11_12_buffer[!clk]) ||(GRF11_13_buffer[clk] != GRF11_13_buffer[!clk]) ||(GRF11_14_buffer[clk] != GRF11_14_buffer[!clk]) ||(GRF11_15_buffer[clk] != GRF11_15_buffer[!clk]) ||(GRF11_16_buffer[clk] != GRF11_16_buffer[!clk]) ||(GRF11_17_buffer[clk] != GRF11_17_buffer[!clk]) ||(GRF11_18_buffer[clk] != GRF11_18_buffer[!clk]) ||(GRF11_19_buffer[clk] != GRF11_19_buffer[!clk]) ||(GRF11_20_buffer[clk] != GRF11_20_buffer[!clk]) ||(GRF11_21_buffer[clk] != GRF11_21_buffer[!clk]) ||(GRF11_22_buffer[clk] != GRF11_22_buffer[!clk]) ||(GRF11_23_buffer[clk] != GRF11_23_buffer[!clk]) ||(GRF11_24_buffer[clk] != GRF11_24_buffer[!clk]) ||(GRF11_25_buffer[clk] != GRF11_25_buffer[!clk]) ||(GRF11_26_buffer[clk] != GRF11_26_buffer[!clk]) ||(GRF11_27_buffer[clk] != GRF11_27_buffer[!clk]) ||(GRF11_28_buffer[clk] != GRF11_28_buffer[!clk]) ||(GRF11_29_buffer[clk] != GRF11_29_buffer[!clk]) ||(GRF11_30_buffer[clk] != GRF11_30_buffer[!clk]) ||(GRF11_31_buffer[clk] != GRF11_31_buffer[!clk]) ||(GRF19_0_buffer[clk] != GRF19_0_buffer[!clk]) ||(GRF19_1_buffer[clk] != GRF19_1_buffer[!clk]) ||(GRF19_2_buffer[clk] != GRF19_2_buffer[!clk]) ||(GRF19_3_buffer[clk] != GRF19_3_buffer[!clk]) ||(GRF19_4_buffer[clk] != GRF19_4_buffer[!clk]) ||(GRF19_5_buffer[clk] != GRF19_5_buffer[!clk]) ||(GRF19_6_buffer[clk] != GRF19_6_buffer[!clk]) ||(GRF19_7_buffer[clk] != GRF19_7_buffer[!clk]) ||(GRF19_8_buffer[clk] != GRF19_8_buffer[!clk]) ||(GRF19_9_buffer[clk] != GRF19_9_buffer[!clk]) ||(GRF19_10_buffer[clk] != GRF19_10_buffer[!clk]) ||(GRF19_11_buffer[clk] != GRF19_11_buffer[!clk]) ||(GRF19_12_buffer[clk] != GRF19_12_buffer[!clk]) ||(GRF19_13_buffer[clk] != GRF19_13_buffer[!clk]) ||(GRF19_14_buffer[clk] != GRF19_14_buffer[!clk]) ||(GRF19_15_buffer[clk] != GRF19_15_buffer[!clk]) ||(GRF19_16_buffer[clk] != GRF19_16_buffer[!clk]) ||(GRF19_17_buffer[clk] != GRF19_17_buffer[!clk]) ||(GRF19_18_buffer[clk] != GRF19_18_buffer[!clk]) ||(GRF19_19_buffer[clk] != GRF19_19_buffer[!clk]) ||(GRF19_20_buffer[clk] != GRF19_20_buffer[!clk]) ||(GRF19_21_buffer[clk] != GRF19_21_buffer[!clk]) ||(GRF19_22_buffer[clk] != GRF19_22_buffer[!clk]) ||(GRF19_23_buffer[clk] != GRF19_23_buffer[!clk]) ||(GRF19_24_buffer[clk] != GRF19_24_buffer[!clk]) ||(GRF19_25_buffer[clk] != GRF19_25_buffer[!clk]) ||(GRF19_26_buffer[clk] != GRF19_26_buffer[!clk]) ||(GRF19_27_buffer[clk] != GRF19_27_buffer[!clk]) ||(GRF19_28_buffer[clk] != GRF19_28_buffer[!clk]) ||(GRF19_29_buffer[clk] != GRF19_29_buffer[!clk]) ||(GRF19_30_buffer[clk] != GRF19_30_buffer[!clk]) ||(GRF19_31_buffer[clk] != GRF19_31_buffer[!clk]) ||(GRF27_0_buffer[clk] != GRF27_0_buffer[!clk]) ||(GRF27_1_buffer[clk] != GRF27_1_buffer[!clk]) ||(GRF27_2_buffer[clk] != GRF27_2_buffer[!clk]) ||(GRF27_3_buffer[clk] != GRF27_3_buffer[!clk]) ||(GRF27_4_buffer[clk] != GRF27_4_buffer[!clk]) ||(GRF27_5_buffer[clk] != GRF27_5_buffer[!clk]) ||(GRF27_6_buffer[clk] != GRF27_6_buffer[!clk]) ||(GRF27_7_buffer[clk] != GRF27_7_buffer[!clk]) ||(GRF27_8_buffer[clk] != GRF27_8_buffer[!clk]) ||(GRF27_9_buffer[clk] != GRF27_9_buffer[!clk]) ||(GRF27_10_buffer[clk] != GRF27_10_buffer[!clk]) ||(GRF27_11_buffer[clk] != GRF27_11_buffer[!clk]) ||(GRF27_12_buffer[clk] != GRF27_12_buffer[!clk]) ||(GRF27_13_buffer[clk] != GRF27_13_buffer[!clk]) ||(GRF27_14_buffer[clk] != GRF27_14_buffer[!clk]) ||(GRF27_15_buffer[clk] != GRF27_15_buffer[!clk]) ||(GRF27_16_buffer[clk] != GRF27_16_buffer[!clk]) ||(GRF27_17_buffer[clk] != GRF27_17_buffer[!clk]) ||(GRF27_18_buffer[clk] != GRF27_18_buffer[!clk]) ||(GRF27_19_buffer[clk] != GRF27_19_buffer[!clk]) ||(GRF27_20_buffer[clk] != GRF27_20_buffer[!clk]) ||(GRF27_21_buffer[clk] != GRF27_21_buffer[!clk]) ||(GRF27_22_buffer[clk] != GRF27_22_buffer[!clk]) ||(GRF27_23_buffer[clk] != GRF27_23_buffer[!clk]) ||(GRF27_24_buffer[clk] != GRF27_24_buffer[!clk]) ||(GRF27_25_buffer[clk] != GRF27_25_buffer[!clk]) ||(GRF27_26_buffer[clk] != GRF27_26_buffer[!clk]) ||(GRF27_27_buffer[clk] != GRF27_27_buffer[!clk]) ||(GRF27_28_buffer[clk] != GRF27_28_buffer[!clk]) ||(GRF27_29_buffer[clk] != GRF27_29_buffer[!clk]) ||(GRF27_30_buffer[clk] != GRF27_30_buffer[!clk]) ||(GRF27_31_buffer[clk] != GRF27_31_buffer[!clk]) ||(GRF35_0_buffer[clk] != GRF35_0_buffer[!clk]) ||(GRF35_1_buffer[clk] != GRF35_1_buffer[!clk]) ||(GRF35_2_buffer[clk] != GRF35_2_buffer[!clk]) ||(GRF35_3_buffer[clk] != GRF35_3_buffer[!clk]) ||(GRF35_4_buffer[clk] != GRF35_4_buffer[!clk]) ||(GRF35_5_buffer[clk] != GRF35_5_buffer[!clk]) ||(GRF35_6_buffer[clk] != GRF35_6_buffer[!clk]) ||(GRF35_7_buffer[clk] != GRF35_7_buffer[!clk]) ||(GRF35_8_buffer[clk] != GRF35_8_buffer[!clk]) ||(GRF35_9_buffer[clk] != GRF35_9_buffer[!clk]) ||(GRF35_10_buffer[clk] != GRF35_10_buffer[!clk]) ||(GRF35_11_buffer[clk] != GRF35_11_buffer[!clk]) ||(GRF35_12_buffer[clk] != GRF35_12_buffer[!clk]) ||(GRF35_13_buffer[clk] != GRF35_13_buffer[!clk]) ||(GRF35_14_buffer[clk] != GRF35_14_buffer[!clk]) ||(GRF35_15_buffer[clk] != GRF35_15_buffer[!clk]) ||(GRF35_16_buffer[clk] != GRF35_16_buffer[!clk]) ||(GRF35_17_buffer[clk] != GRF35_17_buffer[!clk]) ||(GRF35_18_buffer[clk] != GRF35_18_buffer[!clk]) ||(GRF35_19_buffer[clk] != GRF35_19_buffer[!clk]) ||(GRF35_20_buffer[clk] != GRF35_20_buffer[!clk]) ||(GRF35_21_buffer[clk] != GRF35_21_buffer[!clk]) ||(GRF35_22_buffer[clk] != GRF35_22_buffer[!clk]) ||(GRF35_23_buffer[clk] != GRF35_23_buffer[!clk]) ||(GRF35_24_buffer[clk] != GRF35_24_buffer[!clk]) ||(GRF35_25_buffer[clk] != GRF35_25_buffer[!clk]) ||(GRF35_26_buffer[clk] != GRF35_26_buffer[!clk]) ||(GRF35_27_buffer[clk] != GRF35_27_buffer[!clk]) ||(GRF35_28_buffer[clk] != GRF35_28_buffer[!clk]) ||(GRF35_29_buffer[clk] != GRF35_29_buffer[!clk]) ||(GRF35_30_buffer[clk] != GRF35_30_buffer[!clk]) ||(GRF35_31_buffer[clk] != GRF35_31_buffer[!clk]) ||(GRF43_0_buffer[clk] != GRF43_0_buffer[!clk]) ||(GRF43_1_buffer[clk] != GRF43_1_buffer[!clk]) ||(GRF43_2_buffer[clk] != GRF43_2_buffer[!clk]) ||(GRF43_3_buffer[clk] != GRF43_3_buffer[!clk]) ||(GRF43_4_buffer[clk] != GRF43_4_buffer[!clk]) ||(GRF43_5_buffer[clk] != GRF43_5_buffer[!clk]) ||(GRF43_6_buffer[clk] != GRF43_6_buffer[!clk]) ||(GRF43_7_buffer[clk] != GRF43_7_buffer[!clk]) ||(GRF43_8_buffer[clk] != GRF43_8_buffer[!clk]) ||(GRF43_9_buffer[clk] != GRF43_9_buffer[!clk]) ||(GRF43_10_buffer[clk] != GRF43_10_buffer[!clk]) ||(GRF43_11_buffer[clk] != GRF43_11_buffer[!clk]) ||(GRF43_12_buffer[clk] != GRF43_12_buffer[!clk]) ||(GRF43_13_buffer[clk] != GRF43_13_buffer[!clk]) ||(GRF43_14_buffer[clk] != GRF43_14_buffer[!clk]) ||(GRF43_15_buffer[clk] != GRF43_15_buffer[!clk]) ||(GRF43_16_buffer[clk] != GRF43_16_buffer[!clk]) ||(GRF43_17_buffer[clk] != GRF43_17_buffer[!clk]) ||(GRF43_18_buffer[clk] != GRF43_18_buffer[!clk]) ||(GRF43_19_buffer[clk] != GRF43_19_buffer[!clk]) ||(GRF43_20_buffer[clk] != GRF43_20_buffer[!clk]) ||(GRF43_21_buffer[clk] != GRF43_21_buffer[!clk]) ||(GRF43_22_buffer[clk] != GRF43_22_buffer[!clk]) ||(GRF43_23_buffer[clk] != GRF43_23_buffer[!clk]) ||(GRF43_24_buffer[clk] != GRF43_24_buffer[!clk]) ||(GRF43_25_buffer[clk] != GRF43_25_buffer[!clk]) ||(GRF43_26_buffer[clk] != GRF43_26_buffer[!clk]) ||(GRF43_27_buffer[clk] != GRF43_27_buffer[!clk]) ||(GRF43_28_buffer[clk] != GRF43_28_buffer[!clk]) ||(GRF43_29_buffer[clk] != GRF43_29_buffer[!clk]) ||(GRF43_30_buffer[clk] != GRF43_30_buffer[!clk]) ||(GRF43_31_buffer[clk] != GRF43_31_buffer[!clk]) ||(GRF51_0_buffer[clk] != GRF51_0_buffer[!clk]) ||(GRF51_1_buffer[clk] != GRF51_1_buffer[!clk]) ||(GRF51_2_buffer[clk] != GRF51_2_buffer[!clk]) ||(GRF51_3_buffer[clk] != GRF51_3_buffer[!clk]) ||(GRF51_4_buffer[clk] != GRF51_4_buffer[!clk]) ||(GRF51_5_buffer[clk] != GRF51_5_buffer[!clk]) ||(GRF51_6_buffer[clk] != GRF51_6_buffer[!clk]) ||(GRF51_7_buffer[clk] != GRF51_7_buffer[!clk]) ||(GRF51_8_buffer[clk] != GRF51_8_buffer[!clk]) ||(GRF51_9_buffer[clk] != GRF51_9_buffer[!clk]) ||(GRF51_10_buffer[clk] != GRF51_10_buffer[!clk]) ||(GRF51_11_buffer[clk] != GRF51_11_buffer[!clk]) ||(GRF51_12_buffer[clk] != GRF51_12_buffer[!clk]) ||(GRF51_13_buffer[clk] != GRF51_13_buffer[!clk]) ||(GRF51_14_buffer[clk] != GRF51_14_buffer[!clk]) ||(GRF51_15_buffer[clk] != GRF51_15_buffer[!clk]) ||(GRF51_16_buffer[clk] != GRF51_16_buffer[!clk]) ||(GRF51_17_buffer[clk] != GRF51_17_buffer[!clk]) ||(GRF51_18_buffer[clk] != GRF51_18_buffer[!clk]) ||(GRF51_19_buffer[clk] != GRF51_19_buffer[!clk]) ||(GRF51_20_buffer[clk] != GRF51_20_buffer[!clk]) ||(GRF51_21_buffer[clk] != GRF51_21_buffer[!clk]) ||(GRF51_22_buffer[clk] != GRF51_22_buffer[!clk]) ||(GRF51_23_buffer[clk] != GRF51_23_buffer[!clk]) ||(GRF51_24_buffer[clk] != GRF51_24_buffer[!clk]) ||(GRF51_25_buffer[clk] != GRF51_25_buffer[!clk]) ||(GRF51_26_buffer[clk] != GRF51_26_buffer[!clk]) ||(GRF51_27_buffer[clk] != GRF51_27_buffer[!clk]) ||(GRF51_28_buffer[clk] != GRF51_28_buffer[!clk]) ||(GRF51_29_buffer[clk] != GRF51_29_buffer[!clk]) ||(GRF51_30_buffer[clk] != GRF51_30_buffer[!clk]) ||(GRF51_31_buffer[clk] != GRF51_31_buffer[!clk]) ||(GRF59_0_buffer[clk] != GRF59_0_buffer[!clk]) ||(GRF59_1_buffer[clk] != GRF59_1_buffer[!clk]) ||(GRF59_2_buffer[clk] != GRF59_2_buffer[!clk]) ||(GRF59_3_buffer[clk] != GRF59_3_buffer[!clk]) ||(GRF59_4_buffer[clk] != GRF59_4_buffer[!clk]) ||(GRF59_5_buffer[clk] != GRF59_5_buffer[!clk]) ||(GRF59_6_buffer[clk] != GRF59_6_buffer[!clk]) ||(GRF59_7_buffer[clk] != GRF59_7_buffer[!clk]) ||(GRF59_8_buffer[clk] != GRF59_8_buffer[!clk]) ||(GRF59_9_buffer[clk] != GRF59_9_buffer[!clk]) ||(GRF59_10_buffer[clk] != GRF59_10_buffer[!clk]) ||(GRF59_11_buffer[clk] != GRF59_11_buffer[!clk]) ||(GRF59_12_buffer[clk] != GRF59_12_buffer[!clk]) ||(GRF59_13_buffer[clk] != GRF59_13_buffer[!clk]) ||(GRF59_14_buffer[clk] != GRF59_14_buffer[!clk]) ||(GRF59_15_buffer[clk] != GRF59_15_buffer[!clk]) ||(GRF59_16_buffer[clk] != GRF59_16_buffer[!clk]) ||(GRF59_17_buffer[clk] != GRF59_17_buffer[!clk]) ||(GRF59_18_buffer[clk] != GRF59_18_buffer[!clk]) ||(GRF59_19_buffer[clk] != GRF59_19_buffer[!clk]) ||(GRF59_20_buffer[clk] != GRF59_20_buffer[!clk]) ||(GRF59_21_buffer[clk] != GRF59_21_buffer[!clk]) ||(GRF59_22_buffer[clk] != GRF59_22_buffer[!clk]) ||(GRF59_23_buffer[clk] != GRF59_23_buffer[!clk]) ||(GRF59_24_buffer[clk] != GRF59_24_buffer[!clk]) ||(GRF59_25_buffer[clk] != GRF59_25_buffer[!clk]) ||(GRF59_26_buffer[clk] != GRF59_26_buffer[!clk]) ||(GRF59_27_buffer[clk] != GRF59_27_buffer[!clk]) ||(GRF59_28_buffer[clk] != GRF59_28_buffer[!clk]) ||(GRF59_29_buffer[clk] != GRF59_29_buffer[!clk]) ||(GRF59_30_buffer[clk] != GRF59_30_buffer[!clk]) ||(GRF59_31_buffer[clk] != GRF59_31_buffer[!clk]) ) begin
      warp3_sig = 1'b1;
    end else begin
      warp3_sig = 1'b0;
    end

    if ((GRF4_0_buffer[clk] != GRF4_0_buffer[!clk]) ||(GRF4_1_buffer[clk] != GRF4_1_buffer[!clk]) ||(GRF4_2_buffer[clk] != GRF4_2_buffer[!clk]) ||(GRF4_3_buffer[clk] != GRF4_3_buffer[!clk]) ||(GRF4_4_buffer[clk] != GRF4_4_buffer[!clk]) ||(GRF4_5_buffer[clk] != GRF4_5_buffer[!clk]) ||(GRF4_6_buffer[clk] != GRF4_6_buffer[!clk]) ||(GRF4_7_buffer[clk] != GRF4_7_buffer[!clk]) ||(GRF4_8_buffer[clk] != GRF4_8_buffer[!clk]) ||(GRF4_9_buffer[clk] != GRF4_9_buffer[!clk]) ||(GRF4_10_buffer[clk] != GRF4_10_buffer[!clk]) ||(GRF4_11_buffer[clk] != GRF4_11_buffer[!clk]) ||(GRF4_12_buffer[clk] != GRF4_12_buffer[!clk]) ||(GRF4_13_buffer[clk] != GRF4_13_buffer[!clk]) ||(GRF4_14_buffer[clk] != GRF4_14_buffer[!clk]) ||(GRF4_15_buffer[clk] != GRF4_15_buffer[!clk]) ||(GRF4_16_buffer[clk] != GRF4_16_buffer[!clk]) ||(GRF4_17_buffer[clk] != GRF4_17_buffer[!clk]) ||(GRF4_18_buffer[clk] != GRF4_18_buffer[!clk]) ||(GRF4_19_buffer[clk] != GRF4_19_buffer[!clk]) ||(GRF4_20_buffer[clk] != GRF4_20_buffer[!clk]) ||(GRF4_21_buffer[clk] != GRF4_21_buffer[!clk]) ||(GRF4_22_buffer[clk] != GRF4_22_buffer[!clk]) ||(GRF4_23_buffer[clk] != GRF4_23_buffer[!clk]) ||(GRF4_24_buffer[clk] != GRF4_24_buffer[!clk]) ||(GRF4_25_buffer[clk] != GRF4_25_buffer[!clk]) ||(GRF4_26_buffer[clk] != GRF4_26_buffer[!clk]) ||(GRF4_27_buffer[clk] != GRF4_27_buffer[!clk]) ||(GRF4_28_buffer[clk] != GRF4_28_buffer[!clk]) ||(GRF4_29_buffer[clk] != GRF4_29_buffer[!clk]) ||(GRF4_30_buffer[clk] != GRF4_30_buffer[!clk]) ||(GRF4_31_buffer[clk] != GRF4_31_buffer[!clk]) ||(GRF12_0_buffer[clk] != GRF12_0_buffer[!clk]) ||(GRF12_1_buffer[clk] != GRF12_1_buffer[!clk]) ||(GRF12_2_buffer[clk] != GRF12_2_buffer[!clk]) ||(GRF12_3_buffer[clk] != GRF12_3_buffer[!clk]) ||(GRF12_4_buffer[clk] != GRF12_4_buffer[!clk]) ||(GRF12_5_buffer[clk] != GRF12_5_buffer[!clk]) ||(GRF12_6_buffer[clk] != GRF12_6_buffer[!clk]) ||(GRF12_7_buffer[clk] != GRF12_7_buffer[!clk]) ||(GRF12_8_buffer[clk] != GRF12_8_buffer[!clk]) ||(GRF12_9_buffer[clk] != GRF12_9_buffer[!clk]) ||(GRF12_10_buffer[clk] != GRF12_10_buffer[!clk]) ||(GRF12_11_buffer[clk] != GRF12_11_buffer[!clk]) ||(GRF12_12_buffer[clk] != GRF12_12_buffer[!clk]) ||(GRF12_13_buffer[clk] != GRF12_13_buffer[!clk]) ||(GRF12_14_buffer[clk] != GRF12_14_buffer[!clk]) ||(GRF12_15_buffer[clk] != GRF12_15_buffer[!clk]) ||(GRF12_16_buffer[clk] != GRF12_16_buffer[!clk]) ||(GRF12_17_buffer[clk] != GRF12_17_buffer[!clk]) ||(GRF12_18_buffer[clk] != GRF12_18_buffer[!clk]) ||(GRF12_19_buffer[clk] != GRF12_19_buffer[!clk]) ||(GRF12_20_buffer[clk] != GRF12_20_buffer[!clk]) ||(GRF12_21_buffer[clk] != GRF12_21_buffer[!clk]) ||(GRF12_22_buffer[clk] != GRF12_22_buffer[!clk]) ||(GRF12_23_buffer[clk] != GRF12_23_buffer[!clk]) ||(GRF12_24_buffer[clk] != GRF12_24_buffer[!clk]) ||(GRF12_25_buffer[clk] != GRF12_25_buffer[!clk]) ||(GRF12_26_buffer[clk] != GRF12_26_buffer[!clk]) ||(GRF12_27_buffer[clk] != GRF12_27_buffer[!clk]) ||(GRF12_28_buffer[clk] != GRF12_28_buffer[!clk]) ||(GRF12_29_buffer[clk] != GRF12_29_buffer[!clk]) ||(GRF12_30_buffer[clk] != GRF12_30_buffer[!clk]) ||(GRF12_31_buffer[clk] != GRF12_31_buffer[!clk]) ||(GRF20_0_buffer[clk] != GRF20_0_buffer[!clk]) ||(GRF20_1_buffer[clk] != GRF20_1_buffer[!clk]) ||(GRF20_2_buffer[clk] != GRF20_2_buffer[!clk]) ||(GRF20_3_buffer[clk] != GRF20_3_buffer[!clk]) ||(GRF20_4_buffer[clk] != GRF20_4_buffer[!clk]) ||(GRF20_5_buffer[clk] != GRF20_5_buffer[!clk]) ||(GRF20_6_buffer[clk] != GRF20_6_buffer[!clk]) ||(GRF20_7_buffer[clk] != GRF20_7_buffer[!clk]) ||(GRF20_8_buffer[clk] != GRF20_8_buffer[!clk]) ||(GRF20_9_buffer[clk] != GRF20_9_buffer[!clk]) ||(GRF20_10_buffer[clk] != GRF20_10_buffer[!clk]) ||(GRF20_11_buffer[clk] != GRF20_11_buffer[!clk]) ||(GRF20_12_buffer[clk] != GRF20_12_buffer[!clk]) ||(GRF20_13_buffer[clk] != GRF20_13_buffer[!clk]) ||(GRF20_14_buffer[clk] != GRF20_14_buffer[!clk]) ||(GRF20_15_buffer[clk] != GRF20_15_buffer[!clk]) ||(GRF20_16_buffer[clk] != GRF20_16_buffer[!clk]) ||(GRF20_17_buffer[clk] != GRF20_17_buffer[!clk]) ||(GRF20_18_buffer[clk] != GRF20_18_buffer[!clk]) ||(GRF20_19_buffer[clk] != GRF20_19_buffer[!clk]) ||(GRF20_20_buffer[clk] != GRF20_20_buffer[!clk]) ||(GRF20_21_buffer[clk] != GRF20_21_buffer[!clk]) ||(GRF20_22_buffer[clk] != GRF20_22_buffer[!clk]) ||(GRF20_23_buffer[clk] != GRF20_23_buffer[!clk]) ||(GRF20_24_buffer[clk] != GRF20_24_buffer[!clk]) ||(GRF20_25_buffer[clk] != GRF20_25_buffer[!clk]) ||(GRF20_26_buffer[clk] != GRF20_26_buffer[!clk]) ||(GRF20_27_buffer[clk] != GRF20_27_buffer[!clk]) ||(GRF20_28_buffer[clk] != GRF20_28_buffer[!clk]) ||(GRF20_29_buffer[clk] != GRF20_29_buffer[!clk]) ||(GRF20_30_buffer[clk] != GRF20_30_buffer[!clk]) ||(GRF20_31_buffer[clk] != GRF20_31_buffer[!clk]) ||(GRF28_0_buffer[clk] != GRF28_0_buffer[!clk]) ||(GRF28_1_buffer[clk] != GRF28_1_buffer[!clk]) ||(GRF28_2_buffer[clk] != GRF28_2_buffer[!clk]) ||(GRF28_3_buffer[clk] != GRF28_3_buffer[!clk]) ||(GRF28_4_buffer[clk] != GRF28_4_buffer[!clk]) ||(GRF28_5_buffer[clk] != GRF28_5_buffer[!clk]) ||(GRF28_6_buffer[clk] != GRF28_6_buffer[!clk]) ||(GRF28_7_buffer[clk] != GRF28_7_buffer[!clk]) ||(GRF28_8_buffer[clk] != GRF28_8_buffer[!clk]) ||(GRF28_9_buffer[clk] != GRF28_9_buffer[!clk]) ||(GRF28_10_buffer[clk] != GRF28_10_buffer[!clk]) ||(GRF28_11_buffer[clk] != GRF28_11_buffer[!clk]) ||(GRF28_12_buffer[clk] != GRF28_12_buffer[!clk]) ||(GRF28_13_buffer[clk] != GRF28_13_buffer[!clk]) ||(GRF28_14_buffer[clk] != GRF28_14_buffer[!clk]) ||(GRF28_15_buffer[clk] != GRF28_15_buffer[!clk]) ||(GRF28_16_buffer[clk] != GRF28_16_buffer[!clk]) ||(GRF28_17_buffer[clk] != GRF28_17_buffer[!clk]) ||(GRF28_18_buffer[clk] != GRF28_18_buffer[!clk]) ||(GRF28_19_buffer[clk] != GRF28_19_buffer[!clk]) ||(GRF28_20_buffer[clk] != GRF28_20_buffer[!clk]) ||(GRF28_21_buffer[clk] != GRF28_21_buffer[!clk]) ||(GRF28_22_buffer[clk] != GRF28_22_buffer[!clk]) ||(GRF28_23_buffer[clk] != GRF28_23_buffer[!clk]) ||(GRF28_24_buffer[clk] != GRF28_24_buffer[!clk]) ||(GRF28_25_buffer[clk] != GRF28_25_buffer[!clk]) ||(GRF28_26_buffer[clk] != GRF28_26_buffer[!clk]) ||(GRF28_27_buffer[clk] != GRF28_27_buffer[!clk]) ||(GRF28_28_buffer[clk] != GRF28_28_buffer[!clk]) ||(GRF28_29_buffer[clk] != GRF28_29_buffer[!clk]) ||(GRF28_30_buffer[clk] != GRF28_30_buffer[!clk]) ||(GRF28_31_buffer[clk] != GRF28_31_buffer[!clk]) ||(GRF36_0_buffer[clk] != GRF36_0_buffer[!clk]) ||(GRF36_1_buffer[clk] != GRF36_1_buffer[!clk]) ||(GRF36_2_buffer[clk] != GRF36_2_buffer[!clk]) ||(GRF36_3_buffer[clk] != GRF36_3_buffer[!clk]) ||(GRF36_4_buffer[clk] != GRF36_4_buffer[!clk]) ||(GRF36_5_buffer[clk] != GRF36_5_buffer[!clk]) ||(GRF36_6_buffer[clk] != GRF36_6_buffer[!clk]) ||(GRF36_7_buffer[clk] != GRF36_7_buffer[!clk]) ||(GRF36_8_buffer[clk] != GRF36_8_buffer[!clk]) ||(GRF36_9_buffer[clk] != GRF36_9_buffer[!clk]) ||(GRF36_10_buffer[clk] != GRF36_10_buffer[!clk]) ||(GRF36_11_buffer[clk] != GRF36_11_buffer[!clk]) ||(GRF36_12_buffer[clk] != GRF36_12_buffer[!clk]) ||(GRF36_13_buffer[clk] != GRF36_13_buffer[!clk]) ||(GRF36_14_buffer[clk] != GRF36_14_buffer[!clk]) ||(GRF36_15_buffer[clk] != GRF36_15_buffer[!clk]) ||(GRF36_16_buffer[clk] != GRF36_16_buffer[!clk]) ||(GRF36_17_buffer[clk] != GRF36_17_buffer[!clk]) ||(GRF36_18_buffer[clk] != GRF36_18_buffer[!clk]) ||(GRF36_19_buffer[clk] != GRF36_19_buffer[!clk]) ||(GRF36_20_buffer[clk] != GRF36_20_buffer[!clk]) ||(GRF36_21_buffer[clk] != GRF36_21_buffer[!clk]) ||(GRF36_22_buffer[clk] != GRF36_22_buffer[!clk]) ||(GRF36_23_buffer[clk] != GRF36_23_buffer[!clk]) ||(GRF36_24_buffer[clk] != GRF36_24_buffer[!clk]) ||(GRF36_25_buffer[clk] != GRF36_25_buffer[!clk]) ||(GRF36_26_buffer[clk] != GRF36_26_buffer[!clk]) ||(GRF36_27_buffer[clk] != GRF36_27_buffer[!clk]) ||(GRF36_28_buffer[clk] != GRF36_28_buffer[!clk]) ||(GRF36_29_buffer[clk] != GRF36_29_buffer[!clk]) ||(GRF36_30_buffer[clk] != GRF36_30_buffer[!clk]) ||(GRF36_31_buffer[clk] != GRF36_31_buffer[!clk]) ||(GRF44_0_buffer[clk] != GRF44_0_buffer[!clk]) ||(GRF44_1_buffer[clk] != GRF44_1_buffer[!clk]) ||(GRF44_2_buffer[clk] != GRF44_2_buffer[!clk]) ||(GRF44_3_buffer[clk] != GRF44_3_buffer[!clk]) ||(GRF44_4_buffer[clk] != GRF44_4_buffer[!clk]) ||(GRF44_5_buffer[clk] != GRF44_5_buffer[!clk]) ||(GRF44_6_buffer[clk] != GRF44_6_buffer[!clk]) ||(GRF44_7_buffer[clk] != GRF44_7_buffer[!clk]) ||(GRF44_8_buffer[clk] != GRF44_8_buffer[!clk]) ||(GRF44_9_buffer[clk] != GRF44_9_buffer[!clk]) ||(GRF44_10_buffer[clk] != GRF44_10_buffer[!clk]) ||(GRF44_11_buffer[clk] != GRF44_11_buffer[!clk]) ||(GRF44_12_buffer[clk] != GRF44_12_buffer[!clk]) ||(GRF44_13_buffer[clk] != GRF44_13_buffer[!clk]) ||(GRF44_14_buffer[clk] != GRF44_14_buffer[!clk]) ||(GRF44_15_buffer[clk] != GRF44_15_buffer[!clk]) ||(GRF44_16_buffer[clk] != GRF44_16_buffer[!clk]) ||(GRF44_17_buffer[clk] != GRF44_17_buffer[!clk]) ||(GRF44_18_buffer[clk] != GRF44_18_buffer[!clk]) ||(GRF44_19_buffer[clk] != GRF44_19_buffer[!clk]) ||(GRF44_20_buffer[clk] != GRF44_20_buffer[!clk]) ||(GRF44_21_buffer[clk] != GRF44_21_buffer[!clk]) ||(GRF44_22_buffer[clk] != GRF44_22_buffer[!clk]) ||(GRF44_23_buffer[clk] != GRF44_23_buffer[!clk]) ||(GRF44_24_buffer[clk] != GRF44_24_buffer[!clk]) ||(GRF44_25_buffer[clk] != GRF44_25_buffer[!clk]) ||(GRF44_26_buffer[clk] != GRF44_26_buffer[!clk]) ||(GRF44_27_buffer[clk] != GRF44_27_buffer[!clk]) ||(GRF44_28_buffer[clk] != GRF44_28_buffer[!clk]) ||(GRF44_29_buffer[clk] != GRF44_29_buffer[!clk]) ||(GRF44_30_buffer[clk] != GRF44_30_buffer[!clk]) ||(GRF44_31_buffer[clk] != GRF44_31_buffer[!clk]) ||(GRF52_0_buffer[clk] != GRF52_0_buffer[!clk]) ||(GRF52_1_buffer[clk] != GRF52_1_buffer[!clk]) ||(GRF52_2_buffer[clk] != GRF52_2_buffer[!clk]) ||(GRF52_3_buffer[clk] != GRF52_3_buffer[!clk]) ||(GRF52_4_buffer[clk] != GRF52_4_buffer[!clk]) ||(GRF52_5_buffer[clk] != GRF52_5_buffer[!clk]) ||(GRF52_6_buffer[clk] != GRF52_6_buffer[!clk]) ||(GRF52_7_buffer[clk] != GRF52_7_buffer[!clk]) ||(GRF52_8_buffer[clk] != GRF52_8_buffer[!clk]) ||(GRF52_9_buffer[clk] != GRF52_9_buffer[!clk]) ||(GRF52_10_buffer[clk] != GRF52_10_buffer[!clk]) ||(GRF52_11_buffer[clk] != GRF52_11_buffer[!clk]) ||(GRF52_12_buffer[clk] != GRF52_12_buffer[!clk]) ||(GRF52_13_buffer[clk] != GRF52_13_buffer[!clk]) ||(GRF52_14_buffer[clk] != GRF52_14_buffer[!clk]) ||(GRF52_15_buffer[clk] != GRF52_15_buffer[!clk]) ||(GRF52_16_buffer[clk] != GRF52_16_buffer[!clk]) ||(GRF52_17_buffer[clk] != GRF52_17_buffer[!clk]) ||(GRF52_18_buffer[clk] != GRF52_18_buffer[!clk]) ||(GRF52_19_buffer[clk] != GRF52_19_buffer[!clk]) ||(GRF52_20_buffer[clk] != GRF52_20_buffer[!clk]) ||(GRF52_21_buffer[clk] != GRF52_21_buffer[!clk]) ||(GRF52_22_buffer[clk] != GRF52_22_buffer[!clk]) ||(GRF52_23_buffer[clk] != GRF52_23_buffer[!clk]) ||(GRF52_24_buffer[clk] != GRF52_24_buffer[!clk]) ||(GRF52_25_buffer[clk] != GRF52_25_buffer[!clk]) ||(GRF52_26_buffer[clk] != GRF52_26_buffer[!clk]) ||(GRF52_27_buffer[clk] != GRF52_27_buffer[!clk]) ||(GRF52_28_buffer[clk] != GRF52_28_buffer[!clk]) ||(GRF52_29_buffer[clk] != GRF52_29_buffer[!clk]) ||(GRF52_30_buffer[clk] != GRF52_30_buffer[!clk]) ||(GRF52_31_buffer[clk] != GRF52_31_buffer[!clk]) ||(GRF60_0_buffer[clk] != GRF60_0_buffer[!clk]) ||(GRF60_1_buffer[clk] != GRF60_1_buffer[!clk]) ||(GRF60_2_buffer[clk] != GRF60_2_buffer[!clk]) ||(GRF60_3_buffer[clk] != GRF60_3_buffer[!clk]) ||(GRF60_4_buffer[clk] != GRF60_4_buffer[!clk]) ||(GRF60_5_buffer[clk] != GRF60_5_buffer[!clk]) ||(GRF60_6_buffer[clk] != GRF60_6_buffer[!clk]) ||(GRF60_7_buffer[clk] != GRF60_7_buffer[!clk]) ||(GRF60_8_buffer[clk] != GRF60_8_buffer[!clk]) ||(GRF60_9_buffer[clk] != GRF60_9_buffer[!clk]) ||(GRF60_10_buffer[clk] != GRF60_10_buffer[!clk]) ||(GRF60_11_buffer[clk] != GRF60_11_buffer[!clk]) ||(GRF60_12_buffer[clk] != GRF60_12_buffer[!clk]) ||(GRF60_13_buffer[clk] != GRF60_13_buffer[!clk]) ||(GRF60_14_buffer[clk] != GRF60_14_buffer[!clk]) ||(GRF60_15_buffer[clk] != GRF60_15_buffer[!clk]) ||(GRF60_16_buffer[clk] != GRF60_16_buffer[!clk]) ||(GRF60_17_buffer[clk] != GRF60_17_buffer[!clk]) ||(GRF60_18_buffer[clk] != GRF60_18_buffer[!clk]) ||(GRF60_19_buffer[clk] != GRF60_19_buffer[!clk]) ||(GRF60_20_buffer[clk] != GRF60_20_buffer[!clk]) ||(GRF60_21_buffer[clk] != GRF60_21_buffer[!clk]) ||(GRF60_22_buffer[clk] != GRF60_22_buffer[!clk]) ||(GRF60_23_buffer[clk] != GRF60_23_buffer[!clk]) ||(GRF60_24_buffer[clk] != GRF60_24_buffer[!clk]) ||(GRF60_25_buffer[clk] != GRF60_25_buffer[!clk]) ||(GRF60_26_buffer[clk] != GRF60_26_buffer[!clk]) ||(GRF60_27_buffer[clk] != GRF60_27_buffer[!clk]) ||(GRF60_28_buffer[clk] != GRF60_28_buffer[!clk]) ||(GRF60_29_buffer[clk] != GRF60_29_buffer[!clk]) ||(GRF60_30_buffer[clk] != GRF60_30_buffer[!clk]) ||(GRF60_31_buffer[clk] != GRF60_31_buffer[!clk]) ) begin
      warp4_sig = 1'b1;
    end else begin
      warp4_sig = 1'b0;
    end

    if ((GRF5_0_buffer[clk] != GRF5_0_buffer[!clk]) ||(GRF5_1_buffer[clk] != GRF5_1_buffer[!clk]) ||(GRF5_2_buffer[clk] != GRF5_2_buffer[!clk]) ||(GRF5_3_buffer[clk] != GRF5_3_buffer[!clk]) ||(GRF5_4_buffer[clk] != GRF5_4_buffer[!clk]) ||(GRF5_5_buffer[clk] != GRF5_5_buffer[!clk]) ||(GRF5_6_buffer[clk] != GRF5_6_buffer[!clk]) ||(GRF5_7_buffer[clk] != GRF5_7_buffer[!clk]) ||(GRF5_8_buffer[clk] != GRF5_8_buffer[!clk]) ||(GRF5_9_buffer[clk] != GRF5_9_buffer[!clk]) ||(GRF5_10_buffer[clk] != GRF5_10_buffer[!clk]) ||(GRF5_11_buffer[clk] != GRF5_11_buffer[!clk]) ||(GRF5_12_buffer[clk] != GRF5_12_buffer[!clk]) ||(GRF5_13_buffer[clk] != GRF5_13_buffer[!clk]) ||(GRF5_14_buffer[clk] != GRF5_14_buffer[!clk]) ||(GRF5_15_buffer[clk] != GRF5_15_buffer[!clk]) ||(GRF5_16_buffer[clk] != GRF5_16_buffer[!clk]) ||(GRF5_17_buffer[clk] != GRF5_17_buffer[!clk]) ||(GRF5_18_buffer[clk] != GRF5_18_buffer[!clk]) ||(GRF5_19_buffer[clk] != GRF5_19_buffer[!clk]) ||(GRF5_20_buffer[clk] != GRF5_20_buffer[!clk]) ||(GRF5_21_buffer[clk] != GRF5_21_buffer[!clk]) ||(GRF5_22_buffer[clk] != GRF5_22_buffer[!clk]) ||(GRF5_23_buffer[clk] != GRF5_23_buffer[!clk]) ||(GRF5_24_buffer[clk] != GRF5_24_buffer[!clk]) ||(GRF5_25_buffer[clk] != GRF5_25_buffer[!clk]) ||(GRF5_26_buffer[clk] != GRF5_26_buffer[!clk]) ||(GRF5_27_buffer[clk] != GRF5_27_buffer[!clk]) ||(GRF5_28_buffer[clk] != GRF5_28_buffer[!clk]) ||(GRF5_29_buffer[clk] != GRF5_29_buffer[!clk]) ||(GRF5_30_buffer[clk] != GRF5_30_buffer[!clk]) ||(GRF5_31_buffer[clk] != GRF5_31_buffer[!clk]) ||(GRF13_0_buffer[clk] != GRF13_0_buffer[!clk]) ||(GRF13_1_buffer[clk] != GRF13_1_buffer[!clk]) ||(GRF13_2_buffer[clk] != GRF13_2_buffer[!clk]) ||(GRF13_3_buffer[clk] != GRF13_3_buffer[!clk]) ||(GRF13_4_buffer[clk] != GRF13_4_buffer[!clk]) ||(GRF13_5_buffer[clk] != GRF13_5_buffer[!clk]) ||(GRF13_6_buffer[clk] != GRF13_6_buffer[!clk]) ||(GRF13_7_buffer[clk] != GRF13_7_buffer[!clk]) ||(GRF13_8_buffer[clk] != GRF13_8_buffer[!clk]) ||(GRF13_9_buffer[clk] != GRF13_9_buffer[!clk]) ||(GRF13_10_buffer[clk] != GRF13_10_buffer[!clk]) ||(GRF13_11_buffer[clk] != GRF13_11_buffer[!clk]) ||(GRF13_12_buffer[clk] != GRF13_12_buffer[!clk]) ||(GRF13_13_buffer[clk] != GRF13_13_buffer[!clk]) ||(GRF13_14_buffer[clk] != GRF13_14_buffer[!clk]) ||(GRF13_15_buffer[clk] != GRF13_15_buffer[!clk]) ||(GRF13_16_buffer[clk] != GRF13_16_buffer[!clk]) ||(GRF13_17_buffer[clk] != GRF13_17_buffer[!clk]) ||(GRF13_18_buffer[clk] != GRF13_18_buffer[!clk]) ||(GRF13_19_buffer[clk] != GRF13_19_buffer[!clk]) ||(GRF13_20_buffer[clk] != GRF13_20_buffer[!clk]) ||(GRF13_21_buffer[clk] != GRF13_21_buffer[!clk]) ||(GRF13_22_buffer[clk] != GRF13_22_buffer[!clk]) ||(GRF13_23_buffer[clk] != GRF13_23_buffer[!clk]) ||(GRF13_24_buffer[clk] != GRF13_24_buffer[!clk]) ||(GRF13_25_buffer[clk] != GRF13_25_buffer[!clk]) ||(GRF13_26_buffer[clk] != GRF13_26_buffer[!clk]) ||(GRF13_27_buffer[clk] != GRF13_27_buffer[!clk]) ||(GRF13_28_buffer[clk] != GRF13_28_buffer[!clk]) ||(GRF13_29_buffer[clk] != GRF13_29_buffer[!clk]) ||(GRF13_30_buffer[clk] != GRF13_30_buffer[!clk]) ||(GRF13_31_buffer[clk] != GRF13_31_buffer[!clk]) ||(GRF21_0_buffer[clk] != GRF21_0_buffer[!clk]) ||(GRF21_1_buffer[clk] != GRF21_1_buffer[!clk]) ||(GRF21_2_buffer[clk] != GRF21_2_buffer[!clk]) ||(GRF21_3_buffer[clk] != GRF21_3_buffer[!clk]) ||(GRF21_4_buffer[clk] != GRF21_4_buffer[!clk]) ||(GRF21_5_buffer[clk] != GRF21_5_buffer[!clk]) ||(GRF21_6_buffer[clk] != GRF21_6_buffer[!clk]) ||(GRF21_7_buffer[clk] != GRF21_7_buffer[!clk]) ||(GRF21_8_buffer[clk] != GRF21_8_buffer[!clk]) ||(GRF21_9_buffer[clk] != GRF21_9_buffer[!clk]) ||(GRF21_10_buffer[clk] != GRF21_10_buffer[!clk]) ||(GRF21_11_buffer[clk] != GRF21_11_buffer[!clk]) ||(GRF21_12_buffer[clk] != GRF21_12_buffer[!clk]) ||(GRF21_13_buffer[clk] != GRF21_13_buffer[!clk]) ||(GRF21_14_buffer[clk] != GRF21_14_buffer[!clk]) ||(GRF21_15_buffer[clk] != GRF21_15_buffer[!clk]) ||(GRF21_16_buffer[clk] != GRF21_16_buffer[!clk]) ||(GRF21_17_buffer[clk] != GRF21_17_buffer[!clk]) ||(GRF21_18_buffer[clk] != GRF21_18_buffer[!clk]) ||(GRF21_19_buffer[clk] != GRF21_19_buffer[!clk]) ||(GRF21_20_buffer[clk] != GRF21_20_buffer[!clk]) ||(GRF21_21_buffer[clk] != GRF21_21_buffer[!clk]) ||(GRF21_22_buffer[clk] != GRF21_22_buffer[!clk]) ||(GRF21_23_buffer[clk] != GRF21_23_buffer[!clk]) ||(GRF21_24_buffer[clk] != GRF21_24_buffer[!clk]) ||(GRF21_25_buffer[clk] != GRF21_25_buffer[!clk]) ||(GRF21_26_buffer[clk] != GRF21_26_buffer[!clk]) ||(GRF21_27_buffer[clk] != GRF21_27_buffer[!clk]) ||(GRF21_28_buffer[clk] != GRF21_28_buffer[!clk]) ||(GRF21_29_buffer[clk] != GRF21_29_buffer[!clk]) ||(GRF21_30_buffer[clk] != GRF21_30_buffer[!clk]) ||(GRF21_31_buffer[clk] != GRF21_31_buffer[!clk]) ||(GRF29_0_buffer[clk] != GRF29_0_buffer[!clk]) ||(GRF29_1_buffer[clk] != GRF29_1_buffer[!clk]) ||(GRF29_2_buffer[clk] != GRF29_2_buffer[!clk]) ||(GRF29_3_buffer[clk] != GRF29_3_buffer[!clk]) ||(GRF29_4_buffer[clk] != GRF29_4_buffer[!clk]) ||(GRF29_5_buffer[clk] != GRF29_5_buffer[!clk]) ||(GRF29_6_buffer[clk] != GRF29_6_buffer[!clk]) ||(GRF29_7_buffer[clk] != GRF29_7_buffer[!clk]) ||(GRF29_8_buffer[clk] != GRF29_8_buffer[!clk]) ||(GRF29_9_buffer[clk] != GRF29_9_buffer[!clk]) ||(GRF29_10_buffer[clk] != GRF29_10_buffer[!clk]) ||(GRF29_11_buffer[clk] != GRF29_11_buffer[!clk]) ||(GRF29_12_buffer[clk] != GRF29_12_buffer[!clk]) ||(GRF29_13_buffer[clk] != GRF29_13_buffer[!clk]) ||(GRF29_14_buffer[clk] != GRF29_14_buffer[!clk]) ||(GRF29_15_buffer[clk] != GRF29_15_buffer[!clk]) ||(GRF29_16_buffer[clk] != GRF29_16_buffer[!clk]) ||(GRF29_17_buffer[clk] != GRF29_17_buffer[!clk]) ||(GRF29_18_buffer[clk] != GRF29_18_buffer[!clk]) ||(GRF29_19_buffer[clk] != GRF29_19_buffer[!clk]) ||(GRF29_20_buffer[clk] != GRF29_20_buffer[!clk]) ||(GRF29_21_buffer[clk] != GRF29_21_buffer[!clk]) ||(GRF29_22_buffer[clk] != GRF29_22_buffer[!clk]) ||(GRF29_23_buffer[clk] != GRF29_23_buffer[!clk]) ||(GRF29_24_buffer[clk] != GRF29_24_buffer[!clk]) ||(GRF29_25_buffer[clk] != GRF29_25_buffer[!clk]) ||(GRF29_26_buffer[clk] != GRF29_26_buffer[!clk]) ||(GRF29_27_buffer[clk] != GRF29_27_buffer[!clk]) ||(GRF29_28_buffer[clk] != GRF29_28_buffer[!clk]) ||(GRF29_29_buffer[clk] != GRF29_29_buffer[!clk]) ||(GRF29_30_buffer[clk] != GRF29_30_buffer[!clk]) ||(GRF29_31_buffer[clk] != GRF29_31_buffer[!clk]) ||(GRF37_0_buffer[clk] != GRF37_0_buffer[!clk]) ||(GRF37_1_buffer[clk] != GRF37_1_buffer[!clk]) ||(GRF37_2_buffer[clk] != GRF37_2_buffer[!clk]) ||(GRF37_3_buffer[clk] != GRF37_3_buffer[!clk]) ||(GRF37_4_buffer[clk] != GRF37_4_buffer[!clk]) ||(GRF37_5_buffer[clk] != GRF37_5_buffer[!clk]) ||(GRF37_6_buffer[clk] != GRF37_6_buffer[!clk]) ||(GRF37_7_buffer[clk] != GRF37_7_buffer[!clk]) ||(GRF37_8_buffer[clk] != GRF37_8_buffer[!clk]) ||(GRF37_9_buffer[clk] != GRF37_9_buffer[!clk]) ||(GRF37_10_buffer[clk] != GRF37_10_buffer[!clk]) ||(GRF37_11_buffer[clk] != GRF37_11_buffer[!clk]) ||(GRF37_12_buffer[clk] != GRF37_12_buffer[!clk]) ||(GRF37_13_buffer[clk] != GRF37_13_buffer[!clk]) ||(GRF37_14_buffer[clk] != GRF37_14_buffer[!clk]) ||(GRF37_15_buffer[clk] != GRF37_15_buffer[!clk]) ||(GRF37_16_buffer[clk] != GRF37_16_buffer[!clk]) ||(GRF37_17_buffer[clk] != GRF37_17_buffer[!clk]) ||(GRF37_18_buffer[clk] != GRF37_18_buffer[!clk]) ||(GRF37_19_buffer[clk] != GRF37_19_buffer[!clk]) ||(GRF37_20_buffer[clk] != GRF37_20_buffer[!clk]) ||(GRF37_21_buffer[clk] != GRF37_21_buffer[!clk]) ||(GRF37_22_buffer[clk] != GRF37_22_buffer[!clk]) ||(GRF37_23_buffer[clk] != GRF37_23_buffer[!clk]) ||(GRF37_24_buffer[clk] != GRF37_24_buffer[!clk]) ||(GRF37_25_buffer[clk] != GRF37_25_buffer[!clk]) ||(GRF37_26_buffer[clk] != GRF37_26_buffer[!clk]) ||(GRF37_27_buffer[clk] != GRF37_27_buffer[!clk]) ||(GRF37_28_buffer[clk] != GRF37_28_buffer[!clk]) ||(GRF37_29_buffer[clk] != GRF37_29_buffer[!clk]) ||(GRF37_30_buffer[clk] != GRF37_30_buffer[!clk]) ||(GRF37_31_buffer[clk] != GRF37_31_buffer[!clk]) ||(GRF45_0_buffer[clk] != GRF45_0_buffer[!clk]) ||(GRF45_1_buffer[clk] != GRF45_1_buffer[!clk]) ||(GRF45_2_buffer[clk] != GRF45_2_buffer[!clk]) ||(GRF45_3_buffer[clk] != GRF45_3_buffer[!clk]) ||(GRF45_4_buffer[clk] != GRF45_4_buffer[!clk]) ||(GRF45_5_buffer[clk] != GRF45_5_buffer[!clk]) ||(GRF45_6_buffer[clk] != GRF45_6_buffer[!clk]) ||(GRF45_7_buffer[clk] != GRF45_7_buffer[!clk]) ||(GRF45_8_buffer[clk] != GRF45_8_buffer[!clk]) ||(GRF45_9_buffer[clk] != GRF45_9_buffer[!clk]) ||(GRF45_10_buffer[clk] != GRF45_10_buffer[!clk]) ||(GRF45_11_buffer[clk] != GRF45_11_buffer[!clk]) ||(GRF45_12_buffer[clk] != GRF45_12_buffer[!clk]) ||(GRF45_13_buffer[clk] != GRF45_13_buffer[!clk]) ||(GRF45_14_buffer[clk] != GRF45_14_buffer[!clk]) ||(GRF45_15_buffer[clk] != GRF45_15_buffer[!clk]) ||(GRF45_16_buffer[clk] != GRF45_16_buffer[!clk]) ||(GRF45_17_buffer[clk] != GRF45_17_buffer[!clk]) ||(GRF45_18_buffer[clk] != GRF45_18_buffer[!clk]) ||(GRF45_19_buffer[clk] != GRF45_19_buffer[!clk]) ||(GRF45_20_buffer[clk] != GRF45_20_buffer[!clk]) ||(GRF45_21_buffer[clk] != GRF45_21_buffer[!clk]) ||(GRF45_22_buffer[clk] != GRF45_22_buffer[!clk]) ||(GRF45_23_buffer[clk] != GRF45_23_buffer[!clk]) ||(GRF45_24_buffer[clk] != GRF45_24_buffer[!clk]) ||(GRF45_25_buffer[clk] != GRF45_25_buffer[!clk]) ||(GRF45_26_buffer[clk] != GRF45_26_buffer[!clk]) ||(GRF45_27_buffer[clk] != GRF45_27_buffer[!clk]) ||(GRF45_28_buffer[clk] != GRF45_28_buffer[!clk]) ||(GRF45_29_buffer[clk] != GRF45_29_buffer[!clk]) ||(GRF45_30_buffer[clk] != GRF45_30_buffer[!clk]) ||(GRF45_31_buffer[clk] != GRF45_31_buffer[!clk]) ||(GRF53_0_buffer[clk] != GRF53_0_buffer[!clk]) ||(GRF53_1_buffer[clk] != GRF53_1_buffer[!clk]) ||(GRF53_2_buffer[clk] != GRF53_2_buffer[!clk]) ||(GRF53_3_buffer[clk] != GRF53_3_buffer[!clk]) ||(GRF53_4_buffer[clk] != GRF53_4_buffer[!clk]) ||(GRF53_5_buffer[clk] != GRF53_5_buffer[!clk]) ||(GRF53_6_buffer[clk] != GRF53_6_buffer[!clk]) ||(GRF53_7_buffer[clk] != GRF53_7_buffer[!clk]) ||(GRF53_8_buffer[clk] != GRF53_8_buffer[!clk]) ||(GRF53_9_buffer[clk] != GRF53_9_buffer[!clk]) ||(GRF53_10_buffer[clk] != GRF53_10_buffer[!clk]) ||(GRF53_11_buffer[clk] != GRF53_11_buffer[!clk]) ||(GRF53_12_buffer[clk] != GRF53_12_buffer[!clk]) ||(GRF53_13_buffer[clk] != GRF53_13_buffer[!clk]) ||(GRF53_14_buffer[clk] != GRF53_14_buffer[!clk]) ||(GRF53_15_buffer[clk] != GRF53_15_buffer[!clk]) ||(GRF53_16_buffer[clk] != GRF53_16_buffer[!clk]) ||(GRF53_17_buffer[clk] != GRF53_17_buffer[!clk]) ||(GRF53_18_buffer[clk] != GRF53_18_buffer[!clk]) ||(GRF53_19_buffer[clk] != GRF53_19_buffer[!clk]) ||(GRF53_20_buffer[clk] != GRF53_20_buffer[!clk]) ||(GRF53_21_buffer[clk] != GRF53_21_buffer[!clk]) ||(GRF53_22_buffer[clk] != GRF53_22_buffer[!clk]) ||(GRF53_23_buffer[clk] != GRF53_23_buffer[!clk]) ||(GRF53_24_buffer[clk] != GRF53_24_buffer[!clk]) ||(GRF53_25_buffer[clk] != GRF53_25_buffer[!clk]) ||(GRF53_26_buffer[clk] != GRF53_26_buffer[!clk]) ||(GRF53_27_buffer[clk] != GRF53_27_buffer[!clk]) ||(GRF53_28_buffer[clk] != GRF53_28_buffer[!clk]) ||(GRF53_29_buffer[clk] != GRF53_29_buffer[!clk]) ||(GRF53_30_buffer[clk] != GRF53_30_buffer[!clk]) ||(GRF53_31_buffer[clk] != GRF53_31_buffer[!clk]) ||(GRF61_0_buffer[clk] != GRF61_0_buffer[!clk]) ||(GRF61_1_buffer[clk] != GRF61_1_buffer[!clk]) ||(GRF61_2_buffer[clk] != GRF61_2_buffer[!clk]) ||(GRF61_3_buffer[clk] != GRF61_3_buffer[!clk]) ||(GRF61_4_buffer[clk] != GRF61_4_buffer[!clk]) ||(GRF61_5_buffer[clk] != GRF61_5_buffer[!clk]) ||(GRF61_6_buffer[clk] != GRF61_6_buffer[!clk]) ||(GRF61_7_buffer[clk] != GRF61_7_buffer[!clk]) ||(GRF61_8_buffer[clk] != GRF61_8_buffer[!clk]) ||(GRF61_9_buffer[clk] != GRF61_9_buffer[!clk]) ||(GRF61_10_buffer[clk] != GRF61_10_buffer[!clk]) ||(GRF61_11_buffer[clk] != GRF61_11_buffer[!clk]) ||(GRF61_12_buffer[clk] != GRF61_12_buffer[!clk]) ||(GRF61_13_buffer[clk] != GRF61_13_buffer[!clk]) ||(GRF61_14_buffer[clk] != GRF61_14_buffer[!clk]) ||(GRF61_15_buffer[clk] != GRF61_15_buffer[!clk]) ||(GRF61_16_buffer[clk] != GRF61_16_buffer[!clk]) ||(GRF61_17_buffer[clk] != GRF61_17_buffer[!clk]) ||(GRF61_18_buffer[clk] != GRF61_18_buffer[!clk]) ||(GRF61_19_buffer[clk] != GRF61_19_buffer[!clk]) ||(GRF61_20_buffer[clk] != GRF61_20_buffer[!clk]) ||(GRF61_21_buffer[clk] != GRF61_21_buffer[!clk]) ||(GRF61_22_buffer[clk] != GRF61_22_buffer[!clk]) ||(GRF61_23_buffer[clk] != GRF61_23_buffer[!clk]) ||(GRF61_24_buffer[clk] != GRF61_24_buffer[!clk]) ||(GRF61_25_buffer[clk] != GRF61_25_buffer[!clk]) ||(GRF61_26_buffer[clk] != GRF61_26_buffer[!clk]) ||(GRF61_27_buffer[clk] != GRF61_27_buffer[!clk]) ||(GRF61_28_buffer[clk] != GRF61_28_buffer[!clk]) ||(GRF61_29_buffer[clk] != GRF61_29_buffer[!clk]) ||(GRF61_30_buffer[clk] != GRF61_30_buffer[!clk]) ||(GRF61_31_buffer[clk] != GRF61_31_buffer[!clk]) ) begin
      warp5_sig = 1'b1;
    end else begin
      warp5_sig = 1'b0;
    end

    if ((GRF6_0_buffer[clk] != GRF6_0_buffer[!clk]) ||(GRF6_1_buffer[clk] != GRF6_1_buffer[!clk]) ||(GRF6_2_buffer[clk] != GRF6_2_buffer[!clk]) ||(GRF6_3_buffer[clk] != GRF6_3_buffer[!clk]) ||(GRF6_4_buffer[clk] != GRF6_4_buffer[!clk]) ||(GRF6_5_buffer[clk] != GRF6_5_buffer[!clk]) ||(GRF6_6_buffer[clk] != GRF6_6_buffer[!clk]) ||(GRF6_7_buffer[clk] != GRF6_7_buffer[!clk]) ||(GRF6_8_buffer[clk] != GRF6_8_buffer[!clk]) ||(GRF6_9_buffer[clk] != GRF6_9_buffer[!clk]) ||(GRF6_10_buffer[clk] != GRF6_10_buffer[!clk]) ||(GRF6_11_buffer[clk] != GRF6_11_buffer[!clk]) ||(GRF6_12_buffer[clk] != GRF6_12_buffer[!clk]) ||(GRF6_13_buffer[clk] != GRF6_13_buffer[!clk]) ||(GRF6_14_buffer[clk] != GRF6_14_buffer[!clk]) ||(GRF6_15_buffer[clk] != GRF6_15_buffer[!clk]) ||(GRF6_16_buffer[clk] != GRF6_16_buffer[!clk]) ||(GRF6_17_buffer[clk] != GRF6_17_buffer[!clk]) ||(GRF6_18_buffer[clk] != GRF6_18_buffer[!clk]) ||(GRF6_19_buffer[clk] != GRF6_19_buffer[!clk]) ||(GRF6_20_buffer[clk] != GRF6_20_buffer[!clk]) ||(GRF6_21_buffer[clk] != GRF6_21_buffer[!clk]) ||(GRF6_22_buffer[clk] != GRF6_22_buffer[!clk]) ||(GRF6_23_buffer[clk] != GRF6_23_buffer[!clk]) ||(GRF6_24_buffer[clk] != GRF6_24_buffer[!clk]) ||(GRF6_25_buffer[clk] != GRF6_25_buffer[!clk]) ||(GRF6_26_buffer[clk] != GRF6_26_buffer[!clk]) ||(GRF6_27_buffer[clk] != GRF6_27_buffer[!clk]) ||(GRF6_28_buffer[clk] != GRF6_28_buffer[!clk]) ||(GRF6_29_buffer[clk] != GRF6_29_buffer[!clk]) ||(GRF6_30_buffer[clk] != GRF6_30_buffer[!clk]) ||(GRF6_31_buffer[clk] != GRF6_31_buffer[!clk]) ||(GRF14_0_buffer[clk] != GRF14_0_buffer[!clk]) ||(GRF14_1_buffer[clk] != GRF14_1_buffer[!clk]) ||(GRF14_2_buffer[clk] != GRF14_2_buffer[!clk]) ||(GRF14_3_buffer[clk] != GRF14_3_buffer[!clk]) ||(GRF14_4_buffer[clk] != GRF14_4_buffer[!clk]) ||(GRF14_5_buffer[clk] != GRF14_5_buffer[!clk]) ||(GRF14_6_buffer[clk] != GRF14_6_buffer[!clk]) ||(GRF14_7_buffer[clk] != GRF14_7_buffer[!clk]) ||(GRF14_8_buffer[clk] != GRF14_8_buffer[!clk]) ||(GRF14_9_buffer[clk] != GRF14_9_buffer[!clk]) ||(GRF14_10_buffer[clk] != GRF14_10_buffer[!clk]) ||(GRF14_11_buffer[clk] != GRF14_11_buffer[!clk]) ||(GRF14_12_buffer[clk] != GRF14_12_buffer[!clk]) ||(GRF14_13_buffer[clk] != GRF14_13_buffer[!clk]) ||(GRF14_14_buffer[clk] != GRF14_14_buffer[!clk]) ||(GRF14_15_buffer[clk] != GRF14_15_buffer[!clk]) ||(GRF14_16_buffer[clk] != GRF14_16_buffer[!clk]) ||(GRF14_17_buffer[clk] != GRF14_17_buffer[!clk]) ||(GRF14_18_buffer[clk] != GRF14_18_buffer[!clk]) ||(GRF14_19_buffer[clk] != GRF14_19_buffer[!clk]) ||(GRF14_20_buffer[clk] != GRF14_20_buffer[!clk]) ||(GRF14_21_buffer[clk] != GRF14_21_buffer[!clk]) ||(GRF14_22_buffer[clk] != GRF14_22_buffer[!clk]) ||(GRF14_23_buffer[clk] != GRF14_23_buffer[!clk]) ||(GRF14_24_buffer[clk] != GRF14_24_buffer[!clk]) ||(GRF14_25_buffer[clk] != GRF14_25_buffer[!clk]) ||(GRF14_26_buffer[clk] != GRF14_26_buffer[!clk]) ||(GRF14_27_buffer[clk] != GRF14_27_buffer[!clk]) ||(GRF14_28_buffer[clk] != GRF14_28_buffer[!clk]) ||(GRF14_29_buffer[clk] != GRF14_29_buffer[!clk]) ||(GRF14_30_buffer[clk] != GRF14_30_buffer[!clk]) ||(GRF14_31_buffer[clk] != GRF14_31_buffer[!clk]) ||(GRF22_0_buffer[clk] != GRF22_0_buffer[!clk]) ||(GRF22_1_buffer[clk] != GRF22_1_buffer[!clk]) ||(GRF22_2_buffer[clk] != GRF22_2_buffer[!clk]) ||(GRF22_3_buffer[clk] != GRF22_3_buffer[!clk]) ||(GRF22_4_buffer[clk] != GRF22_4_buffer[!clk]) ||(GRF22_5_buffer[clk] != GRF22_5_buffer[!clk]) ||(GRF22_6_buffer[clk] != GRF22_6_buffer[!clk]) ||(GRF22_7_buffer[clk] != GRF22_7_buffer[!clk]) ||(GRF22_8_buffer[clk] != GRF22_8_buffer[!clk]) ||(GRF22_9_buffer[clk] != GRF22_9_buffer[!clk]) ||(GRF22_10_buffer[clk] != GRF22_10_buffer[!clk]) ||(GRF22_11_buffer[clk] != GRF22_11_buffer[!clk]) ||(GRF22_12_buffer[clk] != GRF22_12_buffer[!clk]) ||(GRF22_13_buffer[clk] != GRF22_13_buffer[!clk]) ||(GRF22_14_buffer[clk] != GRF22_14_buffer[!clk]) ||(GRF22_15_buffer[clk] != GRF22_15_buffer[!clk]) ||(GRF22_16_buffer[clk] != GRF22_16_buffer[!clk]) ||(GRF22_17_buffer[clk] != GRF22_17_buffer[!clk]) ||(GRF22_18_buffer[clk] != GRF22_18_buffer[!clk]) ||(GRF22_19_buffer[clk] != GRF22_19_buffer[!clk]) ||(GRF22_20_buffer[clk] != GRF22_20_buffer[!clk]) ||(GRF22_21_buffer[clk] != GRF22_21_buffer[!clk]) ||(GRF22_22_buffer[clk] != GRF22_22_buffer[!clk]) ||(GRF22_23_buffer[clk] != GRF22_23_buffer[!clk]) ||(GRF22_24_buffer[clk] != GRF22_24_buffer[!clk]) ||(GRF22_25_buffer[clk] != GRF22_25_buffer[!clk]) ||(GRF22_26_buffer[clk] != GRF22_26_buffer[!clk]) ||(GRF22_27_buffer[clk] != GRF22_27_buffer[!clk]) ||(GRF22_28_buffer[clk] != GRF22_28_buffer[!clk]) ||(GRF22_29_buffer[clk] != GRF22_29_buffer[!clk]) ||(GRF22_30_buffer[clk] != GRF22_30_buffer[!clk]) ||(GRF22_31_buffer[clk] != GRF22_31_buffer[!clk]) ||(GRF30_0_buffer[clk] != GRF30_0_buffer[!clk]) ||(GRF30_1_buffer[clk] != GRF30_1_buffer[!clk]) ||(GRF30_2_buffer[clk] != GRF30_2_buffer[!clk]) ||(GRF30_3_buffer[clk] != GRF30_3_buffer[!clk]) ||(GRF30_4_buffer[clk] != GRF30_4_buffer[!clk]) ||(GRF30_5_buffer[clk] != GRF30_5_buffer[!clk]) ||(GRF30_6_buffer[clk] != GRF30_6_buffer[!clk]) ||(GRF30_7_buffer[clk] != GRF30_7_buffer[!clk]) ||(GRF30_8_buffer[clk] != GRF30_8_buffer[!clk]) ||(GRF30_9_buffer[clk] != GRF30_9_buffer[!clk]) ||(GRF30_10_buffer[clk] != GRF30_10_buffer[!clk]) ||(GRF30_11_buffer[clk] != GRF30_11_buffer[!clk]) ||(GRF30_12_buffer[clk] != GRF30_12_buffer[!clk]) ||(GRF30_13_buffer[clk] != GRF30_13_buffer[!clk]) ||(GRF30_14_buffer[clk] != GRF30_14_buffer[!clk]) ||(GRF30_15_buffer[clk] != GRF30_15_buffer[!clk]) ||(GRF30_16_buffer[clk] != GRF30_16_buffer[!clk]) ||(GRF30_17_buffer[clk] != GRF30_17_buffer[!clk]) ||(GRF30_18_buffer[clk] != GRF30_18_buffer[!clk]) ||(GRF30_19_buffer[clk] != GRF30_19_buffer[!clk]) ||(GRF30_20_buffer[clk] != GRF30_20_buffer[!clk]) ||(GRF30_21_buffer[clk] != GRF30_21_buffer[!clk]) ||(GRF30_22_buffer[clk] != GRF30_22_buffer[!clk]) ||(GRF30_23_buffer[clk] != GRF30_23_buffer[!clk]) ||(GRF30_24_buffer[clk] != GRF30_24_buffer[!clk]) ||(GRF30_25_buffer[clk] != GRF30_25_buffer[!clk]) ||(GRF30_26_buffer[clk] != GRF30_26_buffer[!clk]) ||(GRF30_27_buffer[clk] != GRF30_27_buffer[!clk]) ||(GRF30_28_buffer[clk] != GRF30_28_buffer[!clk]) ||(GRF30_29_buffer[clk] != GRF30_29_buffer[!clk]) ||(GRF30_30_buffer[clk] != GRF30_30_buffer[!clk]) ||(GRF30_31_buffer[clk] != GRF30_31_buffer[!clk]) ||(GRF38_0_buffer[clk] != GRF38_0_buffer[!clk]) ||(GRF38_1_buffer[clk] != GRF38_1_buffer[!clk]) ||(GRF38_2_buffer[clk] != GRF38_2_buffer[!clk]) ||(GRF38_3_buffer[clk] != GRF38_3_buffer[!clk]) ||(GRF38_4_buffer[clk] != GRF38_4_buffer[!clk]) ||(GRF38_5_buffer[clk] != GRF38_5_buffer[!clk]) ||(GRF38_6_buffer[clk] != GRF38_6_buffer[!clk]) ||(GRF38_7_buffer[clk] != GRF38_7_buffer[!clk]) ||(GRF38_8_buffer[clk] != GRF38_8_buffer[!clk]) ||(GRF38_9_buffer[clk] != GRF38_9_buffer[!clk]) ||(GRF38_10_buffer[clk] != GRF38_10_buffer[!clk]) ||(GRF38_11_buffer[clk] != GRF38_11_buffer[!clk]) ||(GRF38_12_buffer[clk] != GRF38_12_buffer[!clk]) ||(GRF38_13_buffer[clk] != GRF38_13_buffer[!clk]) ||(GRF38_14_buffer[clk] != GRF38_14_buffer[!clk]) ||(GRF38_15_buffer[clk] != GRF38_15_buffer[!clk]) ||(GRF38_16_buffer[clk] != GRF38_16_buffer[!clk]) ||(GRF38_17_buffer[clk] != GRF38_17_buffer[!clk]) ||(GRF38_18_buffer[clk] != GRF38_18_buffer[!clk]) ||(GRF38_19_buffer[clk] != GRF38_19_buffer[!clk]) ||(GRF38_20_buffer[clk] != GRF38_20_buffer[!clk]) ||(GRF38_21_buffer[clk] != GRF38_21_buffer[!clk]) ||(GRF38_22_buffer[clk] != GRF38_22_buffer[!clk]) ||(GRF38_23_buffer[clk] != GRF38_23_buffer[!clk]) ||(GRF38_24_buffer[clk] != GRF38_24_buffer[!clk]) ||(GRF38_25_buffer[clk] != GRF38_25_buffer[!clk]) ||(GRF38_26_buffer[clk] != GRF38_26_buffer[!clk]) ||(GRF38_27_buffer[clk] != GRF38_27_buffer[!clk]) ||(GRF38_28_buffer[clk] != GRF38_28_buffer[!clk]) ||(GRF38_29_buffer[clk] != GRF38_29_buffer[!clk]) ||(GRF38_30_buffer[clk] != GRF38_30_buffer[!clk]) ||(GRF38_31_buffer[clk] != GRF38_31_buffer[!clk]) ||(GRF46_0_buffer[clk] != GRF46_0_buffer[!clk]) ||(GRF46_1_buffer[clk] != GRF46_1_buffer[!clk]) ||(GRF46_2_buffer[clk] != GRF46_2_buffer[!clk]) ||(GRF46_3_buffer[clk] != GRF46_3_buffer[!clk]) ||(GRF46_4_buffer[clk] != GRF46_4_buffer[!clk]) ||(GRF46_5_buffer[clk] != GRF46_5_buffer[!clk]) ||(GRF46_6_buffer[clk] != GRF46_6_buffer[!clk]) ||(GRF46_7_buffer[clk] != GRF46_7_buffer[!clk]) ||(GRF46_8_buffer[clk] != GRF46_8_buffer[!clk]) ||(GRF46_9_buffer[clk] != GRF46_9_buffer[!clk]) ||(GRF46_10_buffer[clk] != GRF46_10_buffer[!clk]) ||(GRF46_11_buffer[clk] != GRF46_11_buffer[!clk]) ||(GRF46_12_buffer[clk] != GRF46_12_buffer[!clk]) ||(GRF46_13_buffer[clk] != GRF46_13_buffer[!clk]) ||(GRF46_14_buffer[clk] != GRF46_14_buffer[!clk]) ||(GRF46_15_buffer[clk] != GRF46_15_buffer[!clk]) ||(GRF46_16_buffer[clk] != GRF46_16_buffer[!clk]) ||(GRF46_17_buffer[clk] != GRF46_17_buffer[!clk]) ||(GRF46_18_buffer[clk] != GRF46_18_buffer[!clk]) ||(GRF46_19_buffer[clk] != GRF46_19_buffer[!clk]) ||(GRF46_20_buffer[clk] != GRF46_20_buffer[!clk]) ||(GRF46_21_buffer[clk] != GRF46_21_buffer[!clk]) ||(GRF46_22_buffer[clk] != GRF46_22_buffer[!clk]) ||(GRF46_23_buffer[clk] != GRF46_23_buffer[!clk]) ||(GRF46_24_buffer[clk] != GRF46_24_buffer[!clk]) ||(GRF46_25_buffer[clk] != GRF46_25_buffer[!clk]) ||(GRF46_26_buffer[clk] != GRF46_26_buffer[!clk]) ||(GRF46_27_buffer[clk] != GRF46_27_buffer[!clk]) ||(GRF46_28_buffer[clk] != GRF46_28_buffer[!clk]) ||(GRF46_29_buffer[clk] != GRF46_29_buffer[!clk]) ||(GRF46_30_buffer[clk] != GRF46_30_buffer[!clk]) ||(GRF46_31_buffer[clk] != GRF46_31_buffer[!clk]) ||(GRF54_0_buffer[clk] != GRF54_0_buffer[!clk]) ||(GRF54_1_buffer[clk] != GRF54_1_buffer[!clk]) ||(GRF54_2_buffer[clk] != GRF54_2_buffer[!clk]) ||(GRF54_3_buffer[clk] != GRF54_3_buffer[!clk]) ||(GRF54_4_buffer[clk] != GRF54_4_buffer[!clk]) ||(GRF54_5_buffer[clk] != GRF54_5_buffer[!clk]) ||(GRF54_6_buffer[clk] != GRF54_6_buffer[!clk]) ||(GRF54_7_buffer[clk] != GRF54_7_buffer[!clk]) ||(GRF54_8_buffer[clk] != GRF54_8_buffer[!clk]) ||(GRF54_9_buffer[clk] != GRF54_9_buffer[!clk]) ||(GRF54_10_buffer[clk] != GRF54_10_buffer[!clk]) ||(GRF54_11_buffer[clk] != GRF54_11_buffer[!clk]) ||(GRF54_12_buffer[clk] != GRF54_12_buffer[!clk]) ||(GRF54_13_buffer[clk] != GRF54_13_buffer[!clk]) ||(GRF54_14_buffer[clk] != GRF54_14_buffer[!clk]) ||(GRF54_15_buffer[clk] != GRF54_15_buffer[!clk]) ||(GRF54_16_buffer[clk] != GRF54_16_buffer[!clk]) ||(GRF54_17_buffer[clk] != GRF54_17_buffer[!clk]) ||(GRF54_18_buffer[clk] != GRF54_18_buffer[!clk]) ||(GRF54_19_buffer[clk] != GRF54_19_buffer[!clk]) ||(GRF54_20_buffer[clk] != GRF54_20_buffer[!clk]) ||(GRF54_21_buffer[clk] != GRF54_21_buffer[!clk]) ||(GRF54_22_buffer[clk] != GRF54_22_buffer[!clk]) ||(GRF54_23_buffer[clk] != GRF54_23_buffer[!clk]) ||(GRF54_24_buffer[clk] != GRF54_24_buffer[!clk]) ||(GRF54_25_buffer[clk] != GRF54_25_buffer[!clk]) ||(GRF54_26_buffer[clk] != GRF54_26_buffer[!clk]) ||(GRF54_27_buffer[clk] != GRF54_27_buffer[!clk]) ||(GRF54_28_buffer[clk] != GRF54_28_buffer[!clk]) ||(GRF54_29_buffer[clk] != GRF54_29_buffer[!clk]) ||(GRF54_30_buffer[clk] != GRF54_30_buffer[!clk]) ||(GRF54_31_buffer[clk] != GRF54_31_buffer[!clk]) ||(GRF62_0_buffer[clk] != GRF62_0_buffer[!clk]) ||(GRF62_1_buffer[clk] != GRF62_1_buffer[!clk]) ||(GRF62_2_buffer[clk] != GRF62_2_buffer[!clk]) ||(GRF62_3_buffer[clk] != GRF62_3_buffer[!clk]) ||(GRF62_4_buffer[clk] != GRF62_4_buffer[!clk]) ||(GRF62_5_buffer[clk] != GRF62_5_buffer[!clk]) ||(GRF62_6_buffer[clk] != GRF62_6_buffer[!clk]) ||(GRF62_7_buffer[clk] != GRF62_7_buffer[!clk]) ||(GRF62_8_buffer[clk] != GRF62_8_buffer[!clk]) ||(GRF62_9_buffer[clk] != GRF62_9_buffer[!clk]) ||(GRF62_10_buffer[clk] != GRF62_10_buffer[!clk]) ||(GRF62_11_buffer[clk] != GRF62_11_buffer[!clk]) ||(GRF62_12_buffer[clk] != GRF62_12_buffer[!clk]) ||(GRF62_13_buffer[clk] != GRF62_13_buffer[!clk]) ||(GRF62_14_buffer[clk] != GRF62_14_buffer[!clk]) ||(GRF62_15_buffer[clk] != GRF62_15_buffer[!clk]) ||(GRF62_16_buffer[clk] != GRF62_16_buffer[!clk]) ||(GRF62_17_buffer[clk] != GRF62_17_buffer[!clk]) ||(GRF62_18_buffer[clk] != GRF62_18_buffer[!clk]) ||(GRF62_19_buffer[clk] != GRF62_19_buffer[!clk]) ||(GRF62_20_buffer[clk] != GRF62_20_buffer[!clk]) ||(GRF62_21_buffer[clk] != GRF62_21_buffer[!clk]) ||(GRF62_22_buffer[clk] != GRF62_22_buffer[!clk]) ||(GRF62_23_buffer[clk] != GRF62_23_buffer[!clk]) ||(GRF62_24_buffer[clk] != GRF62_24_buffer[!clk]) ||(GRF62_25_buffer[clk] != GRF62_25_buffer[!clk]) ||(GRF62_26_buffer[clk] != GRF62_26_buffer[!clk]) ||(GRF62_27_buffer[clk] != GRF62_27_buffer[!clk]) ||(GRF62_28_buffer[clk] != GRF62_28_buffer[!clk]) ||(GRF62_29_buffer[clk] != GRF62_29_buffer[!clk]) ||(GRF62_30_buffer[clk] != GRF62_30_buffer[!clk]) ||(GRF62_31_buffer[clk] != GRF62_31_buffer[!clk]) ) begin
      warp6_sig = 1'b1;
    end else begin
      warp6_sig = 1'b0;
    end

    if ((GRF7_0_buffer[clk] != GRF7_0_buffer[!clk]) ||(GRF7_1_buffer[clk] != GRF7_1_buffer[!clk]) ||(GRF7_2_buffer[clk] != GRF7_2_buffer[!clk]) ||(GRF7_3_buffer[clk] != GRF7_3_buffer[!clk]) ||(GRF7_4_buffer[clk] != GRF7_4_buffer[!clk]) ||(GRF7_5_buffer[clk] != GRF7_5_buffer[!clk]) ||(GRF7_6_buffer[clk] != GRF7_6_buffer[!clk]) ||(GRF7_7_buffer[clk] != GRF7_7_buffer[!clk]) ||(GRF7_8_buffer[clk] != GRF7_8_buffer[!clk]) ||(GRF7_9_buffer[clk] != GRF7_9_buffer[!clk]) ||(GRF7_10_buffer[clk] != GRF7_10_buffer[!clk]) ||(GRF7_11_buffer[clk] != GRF7_11_buffer[!clk]) ||(GRF7_12_buffer[clk] != GRF7_12_buffer[!clk]) ||(GRF7_13_buffer[clk] != GRF7_13_buffer[!clk]) ||(GRF7_14_buffer[clk] != GRF7_14_buffer[!clk]) ||(GRF7_15_buffer[clk] != GRF7_15_buffer[!clk]) ||(GRF7_16_buffer[clk] != GRF7_16_buffer[!clk]) ||(GRF7_17_buffer[clk] != GRF7_17_buffer[!clk]) ||(GRF7_18_buffer[clk] != GRF7_18_buffer[!clk]) ||(GRF7_19_buffer[clk] != GRF7_19_buffer[!clk]) ||(GRF7_20_buffer[clk] != GRF7_20_buffer[!clk]) ||(GRF7_21_buffer[clk] != GRF7_21_buffer[!clk]) ||(GRF7_22_buffer[clk] != GRF7_22_buffer[!clk]) ||(GRF7_23_buffer[clk] != GRF7_23_buffer[!clk]) ||(GRF7_24_buffer[clk] != GRF7_24_buffer[!clk]) ||(GRF7_25_buffer[clk] != GRF7_25_buffer[!clk]) ||(GRF7_26_buffer[clk] != GRF7_26_buffer[!clk]) ||(GRF7_27_buffer[clk] != GRF7_27_buffer[!clk]) ||(GRF7_28_buffer[clk] != GRF7_28_buffer[!clk]) ||(GRF7_29_buffer[clk] != GRF7_29_buffer[!clk]) ||(GRF7_30_buffer[clk] != GRF7_30_buffer[!clk]) ||(GRF7_31_buffer[clk] != GRF7_31_buffer[!clk]) ||(GRF15_0_buffer[clk] != GRF15_0_buffer[!clk]) ||(GRF15_1_buffer[clk] != GRF15_1_buffer[!clk]) ||(GRF15_2_buffer[clk] != GRF15_2_buffer[!clk]) ||(GRF15_3_buffer[clk] != GRF15_3_buffer[!clk]) ||(GRF15_4_buffer[clk] != GRF15_4_buffer[!clk]) ||(GRF15_5_buffer[clk] != GRF15_5_buffer[!clk]) ||(GRF15_6_buffer[clk] != GRF15_6_buffer[!clk]) ||(GRF15_7_buffer[clk] != GRF15_7_buffer[!clk]) ||(GRF15_8_buffer[clk] != GRF15_8_buffer[!clk]) ||(GRF15_9_buffer[clk] != GRF15_9_buffer[!clk]) ||(GRF15_10_buffer[clk] != GRF15_10_buffer[!clk]) ||(GRF15_11_buffer[clk] != GRF15_11_buffer[!clk]) ||(GRF15_12_buffer[clk] != GRF15_12_buffer[!clk]) ||(GRF15_13_buffer[clk] != GRF15_13_buffer[!clk]) ||(GRF15_14_buffer[clk] != GRF15_14_buffer[!clk]) ||(GRF15_15_buffer[clk] != GRF15_15_buffer[!clk]) ||(GRF15_16_buffer[clk] != GRF15_16_buffer[!clk]) ||(GRF15_17_buffer[clk] != GRF15_17_buffer[!clk]) ||(GRF15_18_buffer[clk] != GRF15_18_buffer[!clk]) ||(GRF15_19_buffer[clk] != GRF15_19_buffer[!clk]) ||(GRF15_20_buffer[clk] != GRF15_20_buffer[!clk]) ||(GRF15_21_buffer[clk] != GRF15_21_buffer[!clk]) ||(GRF15_22_buffer[clk] != GRF15_22_buffer[!clk]) ||(GRF15_23_buffer[clk] != GRF15_23_buffer[!clk]) ||(GRF15_24_buffer[clk] != GRF15_24_buffer[!clk]) ||(GRF15_25_buffer[clk] != GRF15_25_buffer[!clk]) ||(GRF15_26_buffer[clk] != GRF15_26_buffer[!clk]) ||(GRF15_27_buffer[clk] != GRF15_27_buffer[!clk]) ||(GRF15_28_buffer[clk] != GRF15_28_buffer[!clk]) ||(GRF15_29_buffer[clk] != GRF15_29_buffer[!clk]) ||(GRF15_30_buffer[clk] != GRF15_30_buffer[!clk]) ||(GRF15_31_buffer[clk] != GRF15_31_buffer[!clk]) ||(GRF23_0_buffer[clk] != GRF23_0_buffer[!clk]) ||(GRF23_1_buffer[clk] != GRF23_1_buffer[!clk]) ||(GRF23_2_buffer[clk] != GRF23_2_buffer[!clk]) ||(GRF23_3_buffer[clk] != GRF23_3_buffer[!clk]) ||(GRF23_4_buffer[clk] != GRF23_4_buffer[!clk]) ||(GRF23_5_buffer[clk] != GRF23_5_buffer[!clk]) ||(GRF23_6_buffer[clk] != GRF23_6_buffer[!clk]) ||(GRF23_7_buffer[clk] != GRF23_7_buffer[!clk]) ||(GRF23_8_buffer[clk] != GRF23_8_buffer[!clk]) ||(GRF23_9_buffer[clk] != GRF23_9_buffer[!clk]) ||(GRF23_10_buffer[clk] != GRF23_10_buffer[!clk]) ||(GRF23_11_buffer[clk] != GRF23_11_buffer[!clk]) ||(GRF23_12_buffer[clk] != GRF23_12_buffer[!clk]) ||(GRF23_13_buffer[clk] != GRF23_13_buffer[!clk]) ||(GRF23_14_buffer[clk] != GRF23_14_buffer[!clk]) ||(GRF23_15_buffer[clk] != GRF23_15_buffer[!clk]) ||(GRF23_16_buffer[clk] != GRF23_16_buffer[!clk]) ||(GRF23_17_buffer[clk] != GRF23_17_buffer[!clk]) ||(GRF23_18_buffer[clk] != GRF23_18_buffer[!clk]) ||(GRF23_19_buffer[clk] != GRF23_19_buffer[!clk]) ||(GRF23_20_buffer[clk] != GRF23_20_buffer[!clk]) ||(GRF23_21_buffer[clk] != GRF23_21_buffer[!clk]) ||(GRF23_22_buffer[clk] != GRF23_22_buffer[!clk]) ||(GRF23_23_buffer[clk] != GRF23_23_buffer[!clk]) ||(GRF23_24_buffer[clk] != GRF23_24_buffer[!clk]) ||(GRF23_25_buffer[clk] != GRF23_25_buffer[!clk]) ||(GRF23_26_buffer[clk] != GRF23_26_buffer[!clk]) ||(GRF23_27_buffer[clk] != GRF23_27_buffer[!clk]) ||(GRF23_28_buffer[clk] != GRF23_28_buffer[!clk]) ||(GRF23_29_buffer[clk] != GRF23_29_buffer[!clk]) ||(GRF23_30_buffer[clk] != GRF23_30_buffer[!clk]) ||(GRF23_31_buffer[clk] != GRF23_31_buffer[!clk]) ||(GRF31_0_buffer[clk] != GRF31_0_buffer[!clk]) ||(GRF31_1_buffer[clk] != GRF31_1_buffer[!clk]) ||(GRF31_2_buffer[clk] != GRF31_2_buffer[!clk]) ||(GRF31_3_buffer[clk] != GRF31_3_buffer[!clk]) ||(GRF31_4_buffer[clk] != GRF31_4_buffer[!clk]) ||(GRF31_5_buffer[clk] != GRF31_5_buffer[!clk]) ||(GRF31_6_buffer[clk] != GRF31_6_buffer[!clk]) ||(GRF31_7_buffer[clk] != GRF31_7_buffer[!clk]) ||(GRF31_8_buffer[clk] != GRF31_8_buffer[!clk]) ||(GRF31_9_buffer[clk] != GRF31_9_buffer[!clk]) ||(GRF31_10_buffer[clk] != GRF31_10_buffer[!clk]) ||(GRF31_11_buffer[clk] != GRF31_11_buffer[!clk]) ||(GRF31_12_buffer[clk] != GRF31_12_buffer[!clk]) ||(GRF31_13_buffer[clk] != GRF31_13_buffer[!clk]) ||(GRF31_14_buffer[clk] != GRF31_14_buffer[!clk]) ||(GRF31_15_buffer[clk] != GRF31_15_buffer[!clk]) ||(GRF31_16_buffer[clk] != GRF31_16_buffer[!clk]) ||(GRF31_17_buffer[clk] != GRF31_17_buffer[!clk]) ||(GRF31_18_buffer[clk] != GRF31_18_buffer[!clk]) ||(GRF31_19_buffer[clk] != GRF31_19_buffer[!clk]) ||(GRF31_20_buffer[clk] != GRF31_20_buffer[!clk]) ||(GRF31_21_buffer[clk] != GRF31_21_buffer[!clk]) ||(GRF31_22_buffer[clk] != GRF31_22_buffer[!clk]) ||(GRF31_23_buffer[clk] != GRF31_23_buffer[!clk]) ||(GRF31_24_buffer[clk] != GRF31_24_buffer[!clk]) ||(GRF31_25_buffer[clk] != GRF31_25_buffer[!clk]) ||(GRF31_26_buffer[clk] != GRF31_26_buffer[!clk]) ||(GRF31_27_buffer[clk] != GRF31_27_buffer[!clk]) ||(GRF31_28_buffer[clk] != GRF31_28_buffer[!clk]) ||(GRF31_29_buffer[clk] != GRF31_29_buffer[!clk]) ||(GRF31_30_buffer[clk] != GRF31_30_buffer[!clk]) ||(GRF31_31_buffer[clk] != GRF31_31_buffer[!clk]) ||(GRF39_0_buffer[clk] != GRF39_0_buffer[!clk]) ||(GRF39_1_buffer[clk] != GRF39_1_buffer[!clk]) ||(GRF39_2_buffer[clk] != GRF39_2_buffer[!clk]) ||(GRF39_3_buffer[clk] != GRF39_3_buffer[!clk]) ||(GRF39_4_buffer[clk] != GRF39_4_buffer[!clk]) ||(GRF39_5_buffer[clk] != GRF39_5_buffer[!clk]) ||(GRF39_6_buffer[clk] != GRF39_6_buffer[!clk]) ||(GRF39_7_buffer[clk] != GRF39_7_buffer[!clk]) ||(GRF39_8_buffer[clk] != GRF39_8_buffer[!clk]) ||(GRF39_9_buffer[clk] != GRF39_9_buffer[!clk]) ||(GRF39_10_buffer[clk] != GRF39_10_buffer[!clk]) ||(GRF39_11_buffer[clk] != GRF39_11_buffer[!clk]) ||(GRF39_12_buffer[clk] != GRF39_12_buffer[!clk]) ||(GRF39_13_buffer[clk] != GRF39_13_buffer[!clk]) ||(GRF39_14_buffer[clk] != GRF39_14_buffer[!clk]) ||(GRF39_15_buffer[clk] != GRF39_15_buffer[!clk]) ||(GRF39_16_buffer[clk] != GRF39_16_buffer[!clk]) ||(GRF39_17_buffer[clk] != GRF39_17_buffer[!clk]) ||(GRF39_18_buffer[clk] != GRF39_18_buffer[!clk]) ||(GRF39_19_buffer[clk] != GRF39_19_buffer[!clk]) ||(GRF39_20_buffer[clk] != GRF39_20_buffer[!clk]) ||(GRF39_21_buffer[clk] != GRF39_21_buffer[!clk]) ||(GRF39_22_buffer[clk] != GRF39_22_buffer[!clk]) ||(GRF39_23_buffer[clk] != GRF39_23_buffer[!clk]) ||(GRF39_24_buffer[clk] != GRF39_24_buffer[!clk]) ||(GRF39_25_buffer[clk] != GRF39_25_buffer[!clk]) ||(GRF39_26_buffer[clk] != GRF39_26_buffer[!clk]) ||(GRF39_27_buffer[clk] != GRF39_27_buffer[!clk]) ||(GRF39_28_buffer[clk] != GRF39_28_buffer[!clk]) ||(GRF39_29_buffer[clk] != GRF39_29_buffer[!clk]) ||(GRF39_30_buffer[clk] != GRF39_30_buffer[!clk]) ||(GRF39_31_buffer[clk] != GRF39_31_buffer[!clk]) ||(GRF47_0_buffer[clk] != GRF47_0_buffer[!clk]) ||(GRF47_1_buffer[clk] != GRF47_1_buffer[!clk]) ||(GRF47_2_buffer[clk] != GRF47_2_buffer[!clk]) ||(GRF47_3_buffer[clk] != GRF47_3_buffer[!clk]) ||(GRF47_4_buffer[clk] != GRF47_4_buffer[!clk]) ||(GRF47_5_buffer[clk] != GRF47_5_buffer[!clk]) ||(GRF47_6_buffer[clk] != GRF47_6_buffer[!clk]) ||(GRF47_7_buffer[clk] != GRF47_7_buffer[!clk]) ||(GRF47_8_buffer[clk] != GRF47_8_buffer[!clk]) ||(GRF47_9_buffer[clk] != GRF47_9_buffer[!clk]) ||(GRF47_10_buffer[clk] != GRF47_10_buffer[!clk]) ||(GRF47_11_buffer[clk] != GRF47_11_buffer[!clk]) ||(GRF47_12_buffer[clk] != GRF47_12_buffer[!clk]) ||(GRF47_13_buffer[clk] != GRF47_13_buffer[!clk]) ||(GRF47_14_buffer[clk] != GRF47_14_buffer[!clk]) ||(GRF47_15_buffer[clk] != GRF47_15_buffer[!clk]) ||(GRF47_16_buffer[clk] != GRF47_16_buffer[!clk]) ||(GRF47_17_buffer[clk] != GRF47_17_buffer[!clk]) ||(GRF47_18_buffer[clk] != GRF47_18_buffer[!clk]) ||(GRF47_19_buffer[clk] != GRF47_19_buffer[!clk]) ||(GRF47_20_buffer[clk] != GRF47_20_buffer[!clk]) ||(GRF47_21_buffer[clk] != GRF47_21_buffer[!clk]) ||(GRF47_22_buffer[clk] != GRF47_22_buffer[!clk]) ||(GRF47_23_buffer[clk] != GRF47_23_buffer[!clk]) ||(GRF47_24_buffer[clk] != GRF47_24_buffer[!clk]) ||(GRF47_25_buffer[clk] != GRF47_25_buffer[!clk]) ||(GRF47_26_buffer[clk] != GRF47_26_buffer[!clk]) ||(GRF47_27_buffer[clk] != GRF47_27_buffer[!clk]) ||(GRF47_28_buffer[clk] != GRF47_28_buffer[!clk]) ||(GRF47_29_buffer[clk] != GRF47_29_buffer[!clk]) ||(GRF47_30_buffer[clk] != GRF47_30_buffer[!clk]) ||(GRF47_31_buffer[clk] != GRF47_31_buffer[!clk]) ||(GRF55_0_buffer[clk] != GRF55_0_buffer[!clk]) ||(GRF55_1_buffer[clk] != GRF55_1_buffer[!clk]) ||(GRF55_2_buffer[clk] != GRF55_2_buffer[!clk]) ||(GRF55_3_buffer[clk] != GRF55_3_buffer[!clk]) ||(GRF55_4_buffer[clk] != GRF55_4_buffer[!clk]) ||(GRF55_5_buffer[clk] != GRF55_5_buffer[!clk]) ||(GRF55_6_buffer[clk] != GRF55_6_buffer[!clk]) ||(GRF55_7_buffer[clk] != GRF55_7_buffer[!clk]) ||(GRF55_8_buffer[clk] != GRF55_8_buffer[!clk]) ||(GRF55_9_buffer[clk] != GRF55_9_buffer[!clk]) ||(GRF55_10_buffer[clk] != GRF55_10_buffer[!clk]) ||(GRF55_11_buffer[clk] != GRF55_11_buffer[!clk]) ||(GRF55_12_buffer[clk] != GRF55_12_buffer[!clk]) ||(GRF55_13_buffer[clk] != GRF55_13_buffer[!clk]) ||(GRF55_14_buffer[clk] != GRF55_14_buffer[!clk]) ||(GRF55_15_buffer[clk] != GRF55_15_buffer[!clk]) ||(GRF55_16_buffer[clk] != GRF55_16_buffer[!clk]) ||(GRF55_17_buffer[clk] != GRF55_17_buffer[!clk]) ||(GRF55_18_buffer[clk] != GRF55_18_buffer[!clk]) ||(GRF55_19_buffer[clk] != GRF55_19_buffer[!clk]) ||(GRF55_20_buffer[clk] != GRF55_20_buffer[!clk]) ||(GRF55_21_buffer[clk] != GRF55_21_buffer[!clk]) ||(GRF55_22_buffer[clk] != GRF55_22_buffer[!clk]) ||(GRF55_23_buffer[clk] != GRF55_23_buffer[!clk]) ||(GRF55_24_buffer[clk] != GRF55_24_buffer[!clk]) ||(GRF55_25_buffer[clk] != GRF55_25_buffer[!clk]) ||(GRF55_26_buffer[clk] != GRF55_26_buffer[!clk]) ||(GRF55_27_buffer[clk] != GRF55_27_buffer[!clk]) ||(GRF55_28_buffer[clk] != GRF55_28_buffer[!clk]) ||(GRF55_29_buffer[clk] != GRF55_29_buffer[!clk]) ||(GRF55_30_buffer[clk] != GRF55_30_buffer[!clk]) ||(GRF55_31_buffer[clk] != GRF55_31_buffer[!clk]) ||(GRF63_0_buffer[clk] != GRF63_0_buffer[!clk]) ||(GRF63_1_buffer[clk] != GRF63_1_buffer[!clk]) ||(GRF63_2_buffer[clk] != GRF63_2_buffer[!clk]) ||(GRF63_3_buffer[clk] != GRF63_3_buffer[!clk]) ||(GRF63_4_buffer[clk] != GRF63_4_buffer[!clk]) ||(GRF63_5_buffer[clk] != GRF63_5_buffer[!clk]) ||(GRF63_6_buffer[clk] != GRF63_6_buffer[!clk]) ||(GRF63_7_buffer[clk] != GRF63_7_buffer[!clk]) ||(GRF63_8_buffer[clk] != GRF63_8_buffer[!clk]) ||(GRF63_9_buffer[clk] != GRF63_9_buffer[!clk]) ||(GRF63_10_buffer[clk] != GRF63_10_buffer[!clk]) ||(GRF63_11_buffer[clk] != GRF63_11_buffer[!clk]) ||(GRF63_12_buffer[clk] != GRF63_12_buffer[!clk]) ||(GRF63_13_buffer[clk] != GRF63_13_buffer[!clk]) ||(GRF63_14_buffer[clk] != GRF63_14_buffer[!clk]) ||(GRF63_15_buffer[clk] != GRF63_15_buffer[!clk]) ||(GRF63_16_buffer[clk] != GRF63_16_buffer[!clk]) ||(GRF63_17_buffer[clk] != GRF63_17_buffer[!clk]) ||(GRF63_18_buffer[clk] != GRF63_18_buffer[!clk]) ||(GRF63_19_buffer[clk] != GRF63_19_buffer[!clk]) ||(GRF63_20_buffer[clk] != GRF63_20_buffer[!clk]) ||(GRF63_21_buffer[clk] != GRF63_21_buffer[!clk]) ||(GRF63_22_buffer[clk] != GRF63_22_buffer[!clk]) ||(GRF63_23_buffer[clk] != GRF63_23_buffer[!clk]) ||(GRF63_24_buffer[clk] != GRF63_24_buffer[!clk]) ||(GRF63_25_buffer[clk] != GRF63_25_buffer[!clk]) ||(GRF63_26_buffer[clk] != GRF63_26_buffer[!clk]) ||(GRF63_27_buffer[clk] != GRF63_27_buffer[!clk]) ||(GRF63_28_buffer[clk] != GRF63_28_buffer[!clk]) ||(GRF63_29_buffer[clk] != GRF63_29_buffer[!clk]) ||(GRF63_30_buffer[clk] != GRF63_30_buffer[!clk]) ||(GRF63_31_buffer[clk] != GRF63_31_buffer[!clk]) ) begin
      warp7_sig = 1'b1;
    end else begin
      warp7_sig = 1'b0;
    end

  end

  // Determine if there is a change in any of the register files
  // When there is a change, then print out the statements below

  // Need to add timestamp, PC start, PC finish, all of Warp Data
  // Output Register Changes
  initial begin
    for (i = 0 ; i < 10000 ; i = i + 1) begin
      @ (posedge clk);
      // pick which warp to trace // WARPEDIT
      if ( warp7_sig == 1'b1 ) begin // change warpX_sig to select
        $fwrite(f, " \n=====================================================\n");
        $fwrite(f, "Simulation Time          ---> ", $time);
        $fwrite(f, "\n\n");

        if (GRF0_0_buffer[clk] != GRF0_0_buffer[!clk]) begin
          $fwrite(f, "Register (0,0) Value: %h\n", GRF0_0_buffer[clk]);
        end
        if (GRF0_1_buffer[clk] != GRF0_1_buffer[!clk]) begin
          $fwrite(f, "Register (0,1) Value: %h\n", GRF0_1_buffer[clk]);
        end
        if (GRF0_2_buffer[clk] != GRF0_2_buffer[!clk]) begin
          $fwrite(f, "Register (0,2) Value: %h\n", GRF0_2_buffer[clk]);
        end
        if (GRF0_3_buffer[clk] != GRF0_3_buffer[!clk]) begin
          $fwrite(f, "Register (0,3) Value: %h\n", GRF0_3_buffer[clk]);
        end
        if (GRF0_4_buffer[clk] != GRF0_4_buffer[!clk]) begin
          $fwrite(f, "Register (0,4) Value: %h\n", GRF0_4_buffer[clk]);
        end
        if (GRF0_5_buffer[clk] != GRF0_5_buffer[!clk]) begin
          $fwrite(f, "Register (0,5) Value: %h\n", GRF0_5_buffer[clk]);
        end
        if (GRF0_6_buffer[clk] != GRF0_6_buffer[!clk]) begin
          $fwrite(f, "Register (0,6) Value: %h\n", GRF0_6_buffer[clk]);
        end
        if (GRF0_7_buffer[clk] != GRF0_7_buffer[!clk]) begin
          $fwrite(f, "Register (0,7) Value: %h\n", GRF0_7_buffer[clk]);
        end
        if (GRF0_8_buffer[clk] != GRF0_8_buffer[!clk]) begin
          $fwrite(f, "Register (0,8) Value: %h\n", GRF0_8_buffer[clk]);
        end
        if (GRF0_9_buffer[clk] != GRF0_9_buffer[!clk]) begin
          $fwrite(f, "Register (0,9) Value: %h\n", GRF0_9_buffer[clk]);
        end
        if (GRF0_10_buffer[clk] != GRF0_10_buffer[!clk]) begin
          $fwrite(f, "Register (0,10) Value: %h\n", GRF0_10_buffer[clk]);
        end
        if (GRF0_11_buffer[clk] != GRF0_11_buffer[!clk]) begin
          $fwrite(f, "Register (0,11) Value: %h\n", GRF0_11_buffer[clk]);
        end
        if (GRF0_12_buffer[clk] != GRF0_12_buffer[!clk]) begin
          $fwrite(f, "Register (0,12) Value: %h\n", GRF0_12_buffer[clk]);
        end
        if (GRF0_13_buffer[clk] != GRF0_13_buffer[!clk]) begin
          $fwrite(f, "Register (0,13) Value: %h\n", GRF0_13_buffer[clk]);
        end
        if (GRF0_14_buffer[clk] != GRF0_14_buffer[!clk]) begin
          $fwrite(f, "Register (0,14) Value: %h\n", GRF0_14_buffer[clk]);
        end
        if (GRF0_15_buffer[clk] != GRF0_15_buffer[!clk]) begin
          $fwrite(f, "Register (0,15) Value: %h\n", GRF0_15_buffer[clk]);
        end
        if (GRF0_16_buffer[clk] != GRF0_16_buffer[!clk]) begin
          $fwrite(f, "Register (0,16) Value: %h\n", GRF0_16_buffer[clk]);
        end
        if (GRF0_17_buffer[clk] != GRF0_17_buffer[!clk]) begin
          $fwrite(f, "Register (0,17) Value: %h\n", GRF0_17_buffer[clk]);
        end
        if (GRF0_18_buffer[clk] != GRF0_18_buffer[!clk]) begin
          $fwrite(f, "Register (0,18) Value: %h\n", GRF0_18_buffer[clk]);
        end
        if (GRF0_19_buffer[clk] != GRF0_19_buffer[!clk]) begin
          $fwrite(f, "Register (0,19) Value: %h\n", GRF0_19_buffer[clk]);
        end
        if (GRF0_20_buffer[clk] != GRF0_20_buffer[!clk]) begin
          $fwrite(f, "Register (0,20) Value: %h\n", GRF0_20_buffer[clk]);
        end
        if (GRF0_21_buffer[clk] != GRF0_21_buffer[!clk]) begin
          $fwrite(f, "Register (0,21) Value: %h\n", GRF0_21_buffer[clk]);
        end
        if (GRF0_22_buffer[clk] != GRF0_22_buffer[!clk]) begin
          $fwrite(f, "Register (0,22) Value: %h\n", GRF0_22_buffer[clk]);
        end
        if (GRF0_23_buffer[clk] != GRF0_23_buffer[!clk]) begin
          $fwrite(f, "Register (0,23) Value: %h\n", GRF0_23_buffer[clk]);
        end
        if (GRF0_24_buffer[clk] != GRF0_24_buffer[!clk]) begin
          $fwrite(f, "Register (0,24) Value: %h\n", GRF0_24_buffer[clk]);
        end
        if (GRF0_25_buffer[clk] != GRF0_25_buffer[!clk]) begin
          $fwrite(f, "Register (0,25) Value: %h\n", GRF0_25_buffer[clk]);
        end
        if (GRF0_26_buffer[clk] != GRF0_26_buffer[!clk]) begin
          $fwrite(f, "Register (0,26) Value: %h\n", GRF0_26_buffer[clk]);
        end
        if (GRF0_27_buffer[clk] != GRF0_27_buffer[!clk]) begin
          $fwrite(f, "Register (0,27) Value: %h\n", GRF0_27_buffer[clk]);
        end
        if (GRF0_28_buffer[clk] != GRF0_28_buffer[!clk]) begin
          $fwrite(f, "Register (0,28) Value: %h\n", GRF0_28_buffer[clk]);
        end
        if (GRF0_29_buffer[clk] != GRF0_29_buffer[!clk]) begin
          $fwrite(f, "Register (0,29) Value: %h\n", GRF0_29_buffer[clk]);
        end
        if (GRF0_30_buffer[clk] != GRF0_30_buffer[!clk]) begin
          $fwrite(f, "Register (0,30) Value: %h\n", GRF0_30_buffer[clk]);
        end
        if (GRF0_31_buffer[clk] != GRF0_31_buffer[!clk]) begin
          $fwrite(f, "Register (0,31) Value: %h\n", GRF0_31_buffer[clk]);
        end
        if (GRF1_0_buffer[clk] != GRF1_0_buffer[!clk]) begin
          $fwrite(f, "Register (1,0) Value: %h\n", GRF1_0_buffer[clk]);
        end
        if (GRF1_1_buffer[clk] != GRF1_1_buffer[!clk]) begin
          $fwrite(f, "Register (1,1) Value: %h\n", GRF1_1_buffer[clk]);
        end
        if (GRF1_2_buffer[clk] != GRF1_2_buffer[!clk]) begin
          $fwrite(f, "Register (1,2) Value: %h\n", GRF1_2_buffer[clk]);
        end
        if (GRF1_3_buffer[clk] != GRF1_3_buffer[!clk]) begin
          $fwrite(f, "Register (1,3) Value: %h\n", GRF1_3_buffer[clk]);
        end
        if (GRF1_4_buffer[clk] != GRF1_4_buffer[!clk]) begin
          $fwrite(f, "Register (1,4) Value: %h\n", GRF1_4_buffer[clk]);
        end
        if (GRF1_5_buffer[clk] != GRF1_5_buffer[!clk]) begin
          $fwrite(f, "Register (1,5) Value: %h\n", GRF1_5_buffer[clk]);
        end
        if (GRF1_6_buffer[clk] != GRF1_6_buffer[!clk]) begin
          $fwrite(f, "Register (1,6) Value: %h\n", GRF1_6_buffer[clk]);
        end
        if (GRF1_7_buffer[clk] != GRF1_7_buffer[!clk]) begin
          $fwrite(f, "Register (1,7) Value: %h\n", GRF1_7_buffer[clk]);
        end
        if (GRF1_8_buffer[clk] != GRF1_8_buffer[!clk]) begin
          $fwrite(f, "Register (1,8) Value: %h\n", GRF1_8_buffer[clk]);
        end
        if (GRF1_9_buffer[clk] != GRF1_9_buffer[!clk]) begin
          $fwrite(f, "Register (1,9) Value: %h\n", GRF1_9_buffer[clk]);
        end
        if (GRF1_10_buffer[clk] != GRF1_10_buffer[!clk]) begin
          $fwrite(f, "Register (1,10) Value: %h\n", GRF1_10_buffer[clk]);
        end
        if (GRF1_11_buffer[clk] != GRF1_11_buffer[!clk]) begin
          $fwrite(f, "Register (1,11) Value: %h\n", GRF1_11_buffer[clk]);
        end
        if (GRF1_12_buffer[clk] != GRF1_12_buffer[!clk]) begin
          $fwrite(f, "Register (1,12) Value: %h\n", GRF1_12_buffer[clk]);
        end
        if (GRF1_13_buffer[clk] != GRF1_13_buffer[!clk]) begin
          $fwrite(f, "Register (1,13) Value: %h\n", GRF1_13_buffer[clk]);
        end
        if (GRF1_14_buffer[clk] != GRF1_14_buffer[!clk]) begin
          $fwrite(f, "Register (1,14) Value: %h\n", GRF1_14_buffer[clk]);
        end
        if (GRF1_15_buffer[clk] != GRF1_15_buffer[!clk]) begin
          $fwrite(f, "Register (1,15) Value: %h\n", GRF1_15_buffer[clk]);
        end
        if (GRF1_16_buffer[clk] != GRF1_16_buffer[!clk]) begin
          $fwrite(f, "Register (1,16) Value: %h\n", GRF1_16_buffer[clk]);
        end
        if (GRF1_17_buffer[clk] != GRF1_17_buffer[!clk]) begin
          $fwrite(f, "Register (1,17) Value: %h\n", GRF1_17_buffer[clk]);
        end
        if (GRF1_18_buffer[clk] != GRF1_18_buffer[!clk]) begin
          $fwrite(f, "Register (1,18) Value: %h\n", GRF1_18_buffer[clk]);
        end
        if (GRF1_19_buffer[clk] != GRF1_19_buffer[!clk]) begin
          $fwrite(f, "Register (1,19) Value: %h\n", GRF1_19_buffer[clk]);
        end
        if (GRF1_20_buffer[clk] != GRF1_20_buffer[!clk]) begin
          $fwrite(f, "Register (1,20) Value: %h\n", GRF1_20_buffer[clk]);
        end
        if (GRF1_21_buffer[clk] != GRF1_21_buffer[!clk]) begin
          $fwrite(f, "Register (1,21) Value: %h\n", GRF1_21_buffer[clk]);
        end
        if (GRF1_22_buffer[clk] != GRF1_22_buffer[!clk]) begin
          $fwrite(f, "Register (1,22) Value: %h\n", GRF1_22_buffer[clk]);
        end
        if (GRF1_23_buffer[clk] != GRF1_23_buffer[!clk]) begin
          $fwrite(f, "Register (1,23) Value: %h\n", GRF1_23_buffer[clk]);
        end
        if (GRF1_24_buffer[clk] != GRF1_24_buffer[!clk]) begin
          $fwrite(f, "Register (1,24) Value: %h\n", GRF1_24_buffer[clk]);
        end
        if (GRF1_25_buffer[clk] != GRF1_25_buffer[!clk]) begin
          $fwrite(f, "Register (1,25) Value: %h\n", GRF1_25_buffer[clk]);
        end
        if (GRF1_26_buffer[clk] != GRF1_26_buffer[!clk]) begin
          $fwrite(f, "Register (1,26) Value: %h\n", GRF1_26_buffer[clk]);
        end
        if (GRF1_27_buffer[clk] != GRF1_27_buffer[!clk]) begin
          $fwrite(f, "Register (1,27) Value: %h\n", GRF1_27_buffer[clk]);
        end
        if (GRF1_28_buffer[clk] != GRF1_28_buffer[!clk]) begin
          $fwrite(f, "Register (1,28) Value: %h\n", GRF1_28_buffer[clk]);
        end
        if (GRF1_29_buffer[clk] != GRF1_29_buffer[!clk]) begin
          $fwrite(f, "Register (1,29) Value: %h\n", GRF1_29_buffer[clk]);
        end
        if (GRF1_30_buffer[clk] != GRF1_30_buffer[!clk]) begin
          $fwrite(f, "Register (1,30) Value: %h\n", GRF1_30_buffer[clk]);
        end
        if (GRF1_31_buffer[clk] != GRF1_31_buffer[!clk]) begin
          $fwrite(f, "Register (1,31) Value: %h\n", GRF1_31_buffer[clk]);
        end
        if (GRF2_0_buffer[clk] != GRF2_0_buffer[!clk]) begin
          $fwrite(f, "Register (2,0) Value: %h\n", GRF2_0_buffer[clk]);
        end
        if (GRF2_1_buffer[clk] != GRF2_1_buffer[!clk]) begin
          $fwrite(f, "Register (2,1) Value: %h\n", GRF2_1_buffer[clk]);
        end
        if (GRF2_2_buffer[clk] != GRF2_2_buffer[!clk]) begin
          $fwrite(f, "Register (2,2) Value: %h\n", GRF2_2_buffer[clk]);
        end
        if (GRF2_3_buffer[clk] != GRF2_3_buffer[!clk]) begin
          $fwrite(f, "Register (2,3) Value: %h\n", GRF2_3_buffer[clk]);
        end
        if (GRF2_4_buffer[clk] != GRF2_4_buffer[!clk]) begin
          $fwrite(f, "Register (2,4) Value: %h\n", GRF2_4_buffer[clk]);
        end
        if (GRF2_5_buffer[clk] != GRF2_5_buffer[!clk]) begin
          $fwrite(f, "Register (2,5) Value: %h\n", GRF2_5_buffer[clk]);
        end
        if (GRF2_6_buffer[clk] != GRF2_6_buffer[!clk]) begin
          $fwrite(f, "Register (2,6) Value: %h\n", GRF2_6_buffer[clk]);
        end
        if (GRF2_7_buffer[clk] != GRF2_7_buffer[!clk]) begin
          $fwrite(f, "Register (2,7) Value: %h\n", GRF2_7_buffer[clk]);
        end
        if (GRF2_8_buffer[clk] != GRF2_8_buffer[!clk]) begin
          $fwrite(f, "Register (2,8) Value: %h\n", GRF2_8_buffer[clk]);
        end
        if (GRF2_9_buffer[clk] != GRF2_9_buffer[!clk]) begin
          $fwrite(f, "Register (2,9) Value: %h\n", GRF2_9_buffer[clk]);
        end
        if (GRF2_10_buffer[clk] != GRF2_10_buffer[!clk]) begin
          $fwrite(f, "Register (2,10) Value: %h\n", GRF2_10_buffer[clk]);
        end
        if (GRF2_11_buffer[clk] != GRF2_11_buffer[!clk]) begin
          $fwrite(f, "Register (2,11) Value: %h\n", GRF2_11_buffer[clk]);
        end
        if (GRF2_12_buffer[clk] != GRF2_12_buffer[!clk]) begin
          $fwrite(f, "Register (2,12) Value: %h\n", GRF2_12_buffer[clk]);
        end
        if (GRF2_13_buffer[clk] != GRF2_13_buffer[!clk]) begin
          $fwrite(f, "Register (2,13) Value: %h\n", GRF2_13_buffer[clk]);
        end
        if (GRF2_14_buffer[clk] != GRF2_14_buffer[!clk]) begin
          $fwrite(f, "Register (2,14) Value: %h\n", GRF2_14_buffer[clk]);
        end
        if (GRF2_15_buffer[clk] != GRF2_15_buffer[!clk]) begin
          $fwrite(f, "Register (2,15) Value: %h\n", GRF2_15_buffer[clk]);
        end
        if (GRF2_16_buffer[clk] != GRF2_16_buffer[!clk]) begin
          $fwrite(f, "Register (2,16) Value: %h\n", GRF2_16_buffer[clk]);
        end
        if (GRF2_17_buffer[clk] != GRF2_17_buffer[!clk]) begin
          $fwrite(f, "Register (2,17) Value: %h\n", GRF2_17_buffer[clk]);
        end
        if (GRF2_18_buffer[clk] != GRF2_18_buffer[!clk]) begin
          $fwrite(f, "Register (2,18) Value: %h\n", GRF2_18_buffer[clk]);
        end
        if (GRF2_19_buffer[clk] != GRF2_19_buffer[!clk]) begin
          $fwrite(f, "Register (2,19) Value: %h\n", GRF2_19_buffer[clk]);
        end
        if (GRF2_20_buffer[clk] != GRF2_20_buffer[!clk]) begin
          $fwrite(f, "Register (2,20) Value: %h\n", GRF2_20_buffer[clk]);
        end
        if (GRF2_21_buffer[clk] != GRF2_21_buffer[!clk]) begin
          $fwrite(f, "Register (2,21) Value: %h\n", GRF2_21_buffer[clk]);
        end
        if (GRF2_22_buffer[clk] != GRF2_22_buffer[!clk]) begin
          $fwrite(f, "Register (2,22) Value: %h\n", GRF2_22_buffer[clk]);
        end
        if (GRF2_23_buffer[clk] != GRF2_23_buffer[!clk]) begin
          $fwrite(f, "Register (2,23) Value: %h\n", GRF2_23_buffer[clk]);
        end
        if (GRF2_24_buffer[clk] != GRF2_24_buffer[!clk]) begin
          $fwrite(f, "Register (2,24) Value: %h\n", GRF2_24_buffer[clk]);
        end
        if (GRF2_25_buffer[clk] != GRF2_25_buffer[!clk]) begin
          $fwrite(f, "Register (2,25) Value: %h\n", GRF2_25_buffer[clk]);
        end
        if (GRF2_26_buffer[clk] != GRF2_26_buffer[!clk]) begin
          $fwrite(f, "Register (2,26) Value: %h\n", GRF2_26_buffer[clk]);
        end
        if (GRF2_27_buffer[clk] != GRF2_27_buffer[!clk]) begin
          $fwrite(f, "Register (2,27) Value: %h\n", GRF2_27_buffer[clk]);
        end
        if (GRF2_28_buffer[clk] != GRF2_28_buffer[!clk]) begin
          $fwrite(f, "Register (2,28) Value: %h\n", GRF2_28_buffer[clk]);
        end
        if (GRF2_29_buffer[clk] != GRF2_29_buffer[!clk]) begin
          $fwrite(f, "Register (2,29) Value: %h\n", GRF2_29_buffer[clk]);
        end
        if (GRF2_30_buffer[clk] != GRF2_30_buffer[!clk]) begin
          $fwrite(f, "Register (2,30) Value: %h\n", GRF2_30_buffer[clk]);
        end
        if (GRF2_31_buffer[clk] != GRF2_31_buffer[!clk]) begin
          $fwrite(f, "Register (2,31) Value: %h\n", GRF2_31_buffer[clk]);
        end
        if (GRF3_0_buffer[clk] != GRF3_0_buffer[!clk]) begin
          $fwrite(f, "Register (3,0) Value: %h\n", GRF3_0_buffer[clk]);
        end
        if (GRF3_1_buffer[clk] != GRF3_1_buffer[!clk]) begin
          $fwrite(f, "Register (3,1) Value: %h\n", GRF3_1_buffer[clk]);
        end
        if (GRF3_2_buffer[clk] != GRF3_2_buffer[!clk]) begin
          $fwrite(f, "Register (3,2) Value: %h\n", GRF3_2_buffer[clk]);
        end
        if (GRF3_3_buffer[clk] != GRF3_3_buffer[!clk]) begin
          $fwrite(f, "Register (3,3) Value: %h\n", GRF3_3_buffer[clk]);
        end
        if (GRF3_4_buffer[clk] != GRF3_4_buffer[!clk]) begin
          $fwrite(f, "Register (3,4) Value: %h\n", GRF3_4_buffer[clk]);
        end
        if (GRF3_5_buffer[clk] != GRF3_5_buffer[!clk]) begin
          $fwrite(f, "Register (3,5) Value: %h\n", GRF3_5_buffer[clk]);
        end
        if (GRF3_6_buffer[clk] != GRF3_6_buffer[!clk]) begin
          $fwrite(f, "Register (3,6) Value: %h\n", GRF3_6_buffer[clk]);
        end
        if (GRF3_7_buffer[clk] != GRF3_7_buffer[!clk]) begin
          $fwrite(f, "Register (3,7) Value: %h\n", GRF3_7_buffer[clk]);
        end
        if (GRF3_8_buffer[clk] != GRF3_8_buffer[!clk]) begin
          $fwrite(f, "Register (3,8) Value: %h\n", GRF3_8_buffer[clk]);
        end
        if (GRF3_9_buffer[clk] != GRF3_9_buffer[!clk]) begin
          $fwrite(f, "Register (3,9) Value: %h\n", GRF3_9_buffer[clk]);
        end
        if (GRF3_10_buffer[clk] != GRF3_10_buffer[!clk]) begin
          $fwrite(f, "Register (3,10) Value: %h\n", GRF3_10_buffer[clk]);
        end
        if (GRF3_11_buffer[clk] != GRF3_11_buffer[!clk]) begin
          $fwrite(f, "Register (3,11) Value: %h\n", GRF3_11_buffer[clk]);
        end
        if (GRF3_12_buffer[clk] != GRF3_12_buffer[!clk]) begin
          $fwrite(f, "Register (3,12) Value: %h\n", GRF3_12_buffer[clk]);
        end
        if (GRF3_13_buffer[clk] != GRF3_13_buffer[!clk]) begin
          $fwrite(f, "Register (3,13) Value: %h\n", GRF3_13_buffer[clk]);
        end
        if (GRF3_14_buffer[clk] != GRF3_14_buffer[!clk]) begin
          $fwrite(f, "Register (3,14) Value: %h\n", GRF3_14_buffer[clk]);
        end
        if (GRF3_15_buffer[clk] != GRF3_15_buffer[!clk]) begin
          $fwrite(f, "Register (3,15) Value: %h\n", GRF3_15_buffer[clk]);
        end
        if (GRF3_16_buffer[clk] != GRF3_16_buffer[!clk]) begin
          $fwrite(f, "Register (3,16) Value: %h\n", GRF3_16_buffer[clk]);
        end
        if (GRF3_17_buffer[clk] != GRF3_17_buffer[!clk]) begin
          $fwrite(f, "Register (3,17) Value: %h\n", GRF3_17_buffer[clk]);
        end
        if (GRF3_18_buffer[clk] != GRF3_18_buffer[!clk]) begin
          $fwrite(f, "Register (3,18) Value: %h\n", GRF3_18_buffer[clk]);
        end
        if (GRF3_19_buffer[clk] != GRF3_19_buffer[!clk]) begin
          $fwrite(f, "Register (3,19) Value: %h\n", GRF3_19_buffer[clk]);
        end
        if (GRF3_20_buffer[clk] != GRF3_20_buffer[!clk]) begin
          $fwrite(f, "Register (3,20) Value: %h\n", GRF3_20_buffer[clk]);
        end
        if (GRF3_21_buffer[clk] != GRF3_21_buffer[!clk]) begin
          $fwrite(f, "Register (3,21) Value: %h\n", GRF3_21_buffer[clk]);
        end
        if (GRF3_22_buffer[clk] != GRF3_22_buffer[!clk]) begin
          $fwrite(f, "Register (3,22) Value: %h\n", GRF3_22_buffer[clk]);
        end
        if (GRF3_23_buffer[clk] != GRF3_23_buffer[!clk]) begin
          $fwrite(f, "Register (3,23) Value: %h\n", GRF3_23_buffer[clk]);
        end
        if (GRF3_24_buffer[clk] != GRF3_24_buffer[!clk]) begin
          $fwrite(f, "Register (3,24) Value: %h\n", GRF3_24_buffer[clk]);
        end
        if (GRF3_25_buffer[clk] != GRF3_25_buffer[!clk]) begin
          $fwrite(f, "Register (3,25) Value: %h\n", GRF3_25_buffer[clk]);
        end
        if (GRF3_26_buffer[clk] != GRF3_26_buffer[!clk]) begin
          $fwrite(f, "Register (3,26) Value: %h\n", GRF3_26_buffer[clk]);
        end
        if (GRF3_27_buffer[clk] != GRF3_27_buffer[!clk]) begin
          $fwrite(f, "Register (3,27) Value: %h\n", GRF3_27_buffer[clk]);
        end
        if (GRF3_28_buffer[clk] != GRF3_28_buffer[!clk]) begin
          $fwrite(f, "Register (3,28) Value: %h\n", GRF3_28_buffer[clk]);
        end
        if (GRF3_29_buffer[clk] != GRF3_29_buffer[!clk]) begin
          $fwrite(f, "Register (3,29) Value: %h\n", GRF3_29_buffer[clk]);
        end
        if (GRF3_30_buffer[clk] != GRF3_30_buffer[!clk]) begin
          $fwrite(f, "Register (3,30) Value: %h\n", GRF3_30_buffer[clk]);
        end
        if (GRF3_31_buffer[clk] != GRF3_31_buffer[!clk]) begin
          $fwrite(f, "Register (3,31) Value: %h\n", GRF3_31_buffer[clk]);
        end
        if (GRF4_0_buffer[clk] != GRF4_0_buffer[!clk]) begin
          $fwrite(f, "Register (4,0) Value: %h\n", GRF4_0_buffer[clk]);
        end
        if (GRF4_1_buffer[clk] != GRF4_1_buffer[!clk]) begin
          $fwrite(f, "Register (4,1) Value: %h\n", GRF4_1_buffer[clk]);
        end
        if (GRF4_2_buffer[clk] != GRF4_2_buffer[!clk]) begin
          $fwrite(f, "Register (4,2) Value: %h\n", GRF4_2_buffer[clk]);
        end
        if (GRF4_3_buffer[clk] != GRF4_3_buffer[!clk]) begin
          $fwrite(f, "Register (4,3) Value: %h\n", GRF4_3_buffer[clk]);
        end
        if (GRF4_4_buffer[clk] != GRF4_4_buffer[!clk]) begin
          $fwrite(f, "Register (4,4) Value: %h\n", GRF4_4_buffer[clk]);
        end
        if (GRF4_5_buffer[clk] != GRF4_5_buffer[!clk]) begin
          $fwrite(f, "Register (4,5) Value: %h\n", GRF4_5_buffer[clk]);
        end
        if (GRF4_6_buffer[clk] != GRF4_6_buffer[!clk]) begin
          $fwrite(f, "Register (4,6) Value: %h\n", GRF4_6_buffer[clk]);
        end
        if (GRF4_7_buffer[clk] != GRF4_7_buffer[!clk]) begin
          $fwrite(f, "Register (4,7) Value: %h\n", GRF4_7_buffer[clk]);
        end
        if (GRF4_8_buffer[clk] != GRF4_8_buffer[!clk]) begin
          $fwrite(f, "Register (4,8) Value: %h\n", GRF4_8_buffer[clk]);
        end
        if (GRF4_9_buffer[clk] != GRF4_9_buffer[!clk]) begin
          $fwrite(f, "Register (4,9) Value: %h\n", GRF4_9_buffer[clk]);
        end
        if (GRF4_10_buffer[clk] != GRF4_10_buffer[!clk]) begin
          $fwrite(f, "Register (4,10) Value: %h\n", GRF4_10_buffer[clk]);
        end
        if (GRF4_11_buffer[clk] != GRF4_11_buffer[!clk]) begin
          $fwrite(f, "Register (4,11) Value: %h\n", GRF4_11_buffer[clk]);
        end
        if (GRF4_12_buffer[clk] != GRF4_12_buffer[!clk]) begin
          $fwrite(f, "Register (4,12) Value: %h\n", GRF4_12_buffer[clk]);
        end
        if (GRF4_13_buffer[clk] != GRF4_13_buffer[!clk]) begin
          $fwrite(f, "Register (4,13) Value: %h\n", GRF4_13_buffer[clk]);
        end
        if (GRF4_14_buffer[clk] != GRF4_14_buffer[!clk]) begin
          $fwrite(f, "Register (4,14) Value: %h\n", GRF4_14_buffer[clk]);
        end
        if (GRF4_15_buffer[clk] != GRF4_15_buffer[!clk]) begin
          $fwrite(f, "Register (4,15) Value: %h\n", GRF4_15_buffer[clk]);
        end
        if (GRF4_16_buffer[clk] != GRF4_16_buffer[!clk]) begin
          $fwrite(f, "Register (4,16) Value: %h\n", GRF4_16_buffer[clk]);
        end
        if (GRF4_17_buffer[clk] != GRF4_17_buffer[!clk]) begin
          $fwrite(f, "Register (4,17) Value: %h\n", GRF4_17_buffer[clk]);
        end
        if (GRF4_18_buffer[clk] != GRF4_18_buffer[!clk]) begin
          $fwrite(f, "Register (4,18) Value: %h\n", GRF4_18_buffer[clk]);
        end
        if (GRF4_19_buffer[clk] != GRF4_19_buffer[!clk]) begin
          $fwrite(f, "Register (4,19) Value: %h\n", GRF4_19_buffer[clk]);
        end
        if (GRF4_20_buffer[clk] != GRF4_20_buffer[!clk]) begin
          $fwrite(f, "Register (4,20) Value: %h\n", GRF4_20_buffer[clk]);
        end
        if (GRF4_21_buffer[clk] != GRF4_21_buffer[!clk]) begin
          $fwrite(f, "Register (4,21) Value: %h\n", GRF4_21_buffer[clk]);
        end
        if (GRF4_22_buffer[clk] != GRF4_22_buffer[!clk]) begin
          $fwrite(f, "Register (4,22) Value: %h\n", GRF4_22_buffer[clk]);
        end
        if (GRF4_23_buffer[clk] != GRF4_23_buffer[!clk]) begin
          $fwrite(f, "Register (4,23) Value: %h\n", GRF4_23_buffer[clk]);
        end
        if (GRF4_24_buffer[clk] != GRF4_24_buffer[!clk]) begin
          $fwrite(f, "Register (4,24) Value: %h\n", GRF4_24_buffer[clk]);
        end
        if (GRF4_25_buffer[clk] != GRF4_25_buffer[!clk]) begin
          $fwrite(f, "Register (4,25) Value: %h\n", GRF4_25_buffer[clk]);
        end
        if (GRF4_26_buffer[clk] != GRF4_26_buffer[!clk]) begin
          $fwrite(f, "Register (4,26) Value: %h\n", GRF4_26_buffer[clk]);
        end
        if (GRF4_27_buffer[clk] != GRF4_27_buffer[!clk]) begin
          $fwrite(f, "Register (4,27) Value: %h\n", GRF4_27_buffer[clk]);
        end
        if (GRF4_28_buffer[clk] != GRF4_28_buffer[!clk]) begin
          $fwrite(f, "Register (4,28) Value: %h\n", GRF4_28_buffer[clk]);
        end
        if (GRF4_29_buffer[clk] != GRF4_29_buffer[!clk]) begin
          $fwrite(f, "Register (4,29) Value: %h\n", GRF4_29_buffer[clk]);
        end
        if (GRF4_30_buffer[clk] != GRF4_30_buffer[!clk]) begin
          $fwrite(f, "Register (4,30) Value: %h\n", GRF4_30_buffer[clk]);
        end
        if (GRF4_31_buffer[clk] != GRF4_31_buffer[!clk]) begin
          $fwrite(f, "Register (4,31) Value: %h\n", GRF4_31_buffer[clk]);
        end
        if (GRF5_0_buffer[clk] != GRF5_0_buffer[!clk]) begin
          $fwrite(f, "Register (5,0) Value: %h\n", GRF5_0_buffer[clk]);
        end
        if (GRF5_1_buffer[clk] != GRF5_1_buffer[!clk]) begin
          $fwrite(f, "Register (5,1) Value: %h\n", GRF5_1_buffer[clk]);
        end
        if (GRF5_2_buffer[clk] != GRF5_2_buffer[!clk]) begin
          $fwrite(f, "Register (5,2) Value: %h\n", GRF5_2_buffer[clk]);
        end
        if (GRF5_3_buffer[clk] != GRF5_3_buffer[!clk]) begin
          $fwrite(f, "Register (5,3) Value: %h\n", GRF5_3_buffer[clk]);
        end
        if (GRF5_4_buffer[clk] != GRF5_4_buffer[!clk]) begin
          $fwrite(f, "Register (5,4) Value: %h\n", GRF5_4_buffer[clk]);
        end
        if (GRF5_5_buffer[clk] != GRF5_5_buffer[!clk]) begin
          $fwrite(f, "Register (5,5) Value: %h\n", GRF5_5_buffer[clk]);
        end
        if (GRF5_6_buffer[clk] != GRF5_6_buffer[!clk]) begin
          $fwrite(f, "Register (5,6) Value: %h\n", GRF5_6_buffer[clk]);
        end
        if (GRF5_7_buffer[clk] != GRF5_7_buffer[!clk]) begin
          $fwrite(f, "Register (5,7) Value: %h\n", GRF5_7_buffer[clk]);
        end
        if (GRF5_8_buffer[clk] != GRF5_8_buffer[!clk]) begin
          $fwrite(f, "Register (5,8) Value: %h\n", GRF5_8_buffer[clk]);
        end
        if (GRF5_9_buffer[clk] != GRF5_9_buffer[!clk]) begin
          $fwrite(f, "Register (5,9) Value: %h\n", GRF5_9_buffer[clk]);
        end
        if (GRF5_10_buffer[clk] != GRF5_10_buffer[!clk]) begin
          $fwrite(f, "Register (5,10) Value: %h\n", GRF5_10_buffer[clk]);
        end
        if (GRF5_11_buffer[clk] != GRF5_11_buffer[!clk]) begin
          $fwrite(f, "Register (5,11) Value: %h\n", GRF5_11_buffer[clk]);
        end
        if (GRF5_12_buffer[clk] != GRF5_12_buffer[!clk]) begin
          $fwrite(f, "Register (5,12) Value: %h\n", GRF5_12_buffer[clk]);
        end
        if (GRF5_13_buffer[clk] != GRF5_13_buffer[!clk]) begin
          $fwrite(f, "Register (5,13) Value: %h\n", GRF5_13_buffer[clk]);
        end
        if (GRF5_14_buffer[clk] != GRF5_14_buffer[!clk]) begin
          $fwrite(f, "Register (5,14) Value: %h\n", GRF5_14_buffer[clk]);
        end
        if (GRF5_15_buffer[clk] != GRF5_15_buffer[!clk]) begin
          $fwrite(f, "Register (5,15) Value: %h\n", GRF5_15_buffer[clk]);
        end
        if (GRF5_16_buffer[clk] != GRF5_16_buffer[!clk]) begin
          $fwrite(f, "Register (5,16) Value: %h\n", GRF5_16_buffer[clk]);
        end
        if (GRF5_17_buffer[clk] != GRF5_17_buffer[!clk]) begin
          $fwrite(f, "Register (5,17) Value: %h\n", GRF5_17_buffer[clk]);
        end
        if (GRF5_18_buffer[clk] != GRF5_18_buffer[!clk]) begin
          $fwrite(f, "Register (5,18) Value: %h\n", GRF5_18_buffer[clk]);
        end
        if (GRF5_19_buffer[clk] != GRF5_19_buffer[!clk]) begin
          $fwrite(f, "Register (5,19) Value: %h\n", GRF5_19_buffer[clk]);
        end
        if (GRF5_20_buffer[clk] != GRF5_20_buffer[!clk]) begin
          $fwrite(f, "Register (5,20) Value: %h\n", GRF5_20_buffer[clk]);
        end
        if (GRF5_21_buffer[clk] != GRF5_21_buffer[!clk]) begin
          $fwrite(f, "Register (5,21) Value: %h\n", GRF5_21_buffer[clk]);
        end
        if (GRF5_22_buffer[clk] != GRF5_22_buffer[!clk]) begin
          $fwrite(f, "Register (5,22) Value: %h\n", GRF5_22_buffer[clk]);
        end
        if (GRF5_23_buffer[clk] != GRF5_23_buffer[!clk]) begin
          $fwrite(f, "Register (5,23) Value: %h\n", GRF5_23_buffer[clk]);
        end
        if (GRF5_24_buffer[clk] != GRF5_24_buffer[!clk]) begin
          $fwrite(f, "Register (5,24) Value: %h\n", GRF5_24_buffer[clk]);
        end
        if (GRF5_25_buffer[clk] != GRF5_25_buffer[!clk]) begin
          $fwrite(f, "Register (5,25) Value: %h\n", GRF5_25_buffer[clk]);
        end
        if (GRF5_26_buffer[clk] != GRF5_26_buffer[!clk]) begin
          $fwrite(f, "Register (5,26) Value: %h\n", GRF5_26_buffer[clk]);
        end
        if (GRF5_27_buffer[clk] != GRF5_27_buffer[!clk]) begin
          $fwrite(f, "Register (5,27) Value: %h\n", GRF5_27_buffer[clk]);
        end
        if (GRF5_28_buffer[clk] != GRF5_28_buffer[!clk]) begin
          $fwrite(f, "Register (5,28) Value: %h\n", GRF5_28_buffer[clk]);
        end
        if (GRF5_29_buffer[clk] != GRF5_29_buffer[!clk]) begin
          $fwrite(f, "Register (5,29) Value: %h\n", GRF5_29_buffer[clk]);
        end
        if (GRF5_30_buffer[clk] != GRF5_30_buffer[!clk]) begin
          $fwrite(f, "Register (5,30) Value: %h\n", GRF5_30_buffer[clk]);
        end
        if (GRF5_31_buffer[clk] != GRF5_31_buffer[!clk]) begin
          $fwrite(f, "Register (5,31) Value: %h\n", GRF5_31_buffer[clk]);
        end
        if (GRF6_0_buffer[clk] != GRF6_0_buffer[!clk]) begin
          $fwrite(f, "Register (6,0) Value: %h\n", GRF6_0_buffer[clk]);
        end
        if (GRF6_1_buffer[clk] != GRF6_1_buffer[!clk]) begin
          $fwrite(f, "Register (6,1) Value: %h\n", GRF6_1_buffer[clk]);
        end
        if (GRF6_2_buffer[clk] != GRF6_2_buffer[!clk]) begin
          $fwrite(f, "Register (6,2) Value: %h\n", GRF6_2_buffer[clk]);
        end
        if (GRF6_3_buffer[clk] != GRF6_3_buffer[!clk]) begin
          $fwrite(f, "Register (6,3) Value: %h\n", GRF6_3_buffer[clk]);
        end
        if (GRF6_4_buffer[clk] != GRF6_4_buffer[!clk]) begin
          $fwrite(f, "Register (6,4) Value: %h\n", GRF6_4_buffer[clk]);
        end
        if (GRF6_5_buffer[clk] != GRF6_5_buffer[!clk]) begin
          $fwrite(f, "Register (6,5) Value: %h\n", GRF6_5_buffer[clk]);
        end
        if (GRF6_6_buffer[clk] != GRF6_6_buffer[!clk]) begin
          $fwrite(f, "Register (6,6) Value: %h\n", GRF6_6_buffer[clk]);
        end
        if (GRF6_7_buffer[clk] != GRF6_7_buffer[!clk]) begin
          $fwrite(f, "Register (6,7) Value: %h\n", GRF6_7_buffer[clk]);
        end
        if (GRF6_8_buffer[clk] != GRF6_8_buffer[!clk]) begin
          $fwrite(f, "Register (6,8) Value: %h\n", GRF6_8_buffer[clk]);
        end
        if (GRF6_9_buffer[clk] != GRF6_9_buffer[!clk]) begin
          $fwrite(f, "Register (6,9) Value: %h\n", GRF6_9_buffer[clk]);
        end
        if (GRF6_10_buffer[clk] != GRF6_10_buffer[!clk]) begin
          $fwrite(f, "Register (6,10) Value: %h\n", GRF6_10_buffer[clk]);
        end
        if (GRF6_11_buffer[clk] != GRF6_11_buffer[!clk]) begin
          $fwrite(f, "Register (6,11) Value: %h\n", GRF6_11_buffer[clk]);
        end
        if (GRF6_12_buffer[clk] != GRF6_12_buffer[!clk]) begin
          $fwrite(f, "Register (6,12) Value: %h\n", GRF6_12_buffer[clk]);
        end
        if (GRF6_13_buffer[clk] != GRF6_13_buffer[!clk]) begin
          $fwrite(f, "Register (6,13) Value: %h\n", GRF6_13_buffer[clk]);
        end
        if (GRF6_14_buffer[clk] != GRF6_14_buffer[!clk]) begin
          $fwrite(f, "Register (6,14) Value: %h\n", GRF6_14_buffer[clk]);
        end
        if (GRF6_15_buffer[clk] != GRF6_15_buffer[!clk]) begin
          $fwrite(f, "Register (6,15) Value: %h\n", GRF6_15_buffer[clk]);
        end
        if (GRF6_16_buffer[clk] != GRF6_16_buffer[!clk]) begin
          $fwrite(f, "Register (6,16) Value: %h\n", GRF6_16_buffer[clk]);
        end
        if (GRF6_17_buffer[clk] != GRF6_17_buffer[!clk]) begin
          $fwrite(f, "Register (6,17) Value: %h\n", GRF6_17_buffer[clk]);
        end
        if (GRF6_18_buffer[clk] != GRF6_18_buffer[!clk]) begin
          $fwrite(f, "Register (6,18) Value: %h\n", GRF6_18_buffer[clk]);
        end
        if (GRF6_19_buffer[clk] != GRF6_19_buffer[!clk]) begin
          $fwrite(f, "Register (6,19) Value: %h\n", GRF6_19_buffer[clk]);
        end
        if (GRF6_20_buffer[clk] != GRF6_20_buffer[!clk]) begin
          $fwrite(f, "Register (6,20) Value: %h\n", GRF6_20_buffer[clk]);
        end
        if (GRF6_21_buffer[clk] != GRF6_21_buffer[!clk]) begin
          $fwrite(f, "Register (6,21) Value: %h\n", GRF6_21_buffer[clk]);
        end
        if (GRF6_22_buffer[clk] != GRF6_22_buffer[!clk]) begin
          $fwrite(f, "Register (6,22) Value: %h\n", GRF6_22_buffer[clk]);
        end
        if (GRF6_23_buffer[clk] != GRF6_23_buffer[!clk]) begin
          $fwrite(f, "Register (6,23) Value: %h\n", GRF6_23_buffer[clk]);
        end
        if (GRF6_24_buffer[clk] != GRF6_24_buffer[!clk]) begin
          $fwrite(f, "Register (6,24) Value: %h\n", GRF6_24_buffer[clk]);
        end
        if (GRF6_25_buffer[clk] != GRF6_25_buffer[!clk]) begin
          $fwrite(f, "Register (6,25) Value: %h\n", GRF6_25_buffer[clk]);
        end
        if (GRF6_26_buffer[clk] != GRF6_26_buffer[!clk]) begin
          $fwrite(f, "Register (6,26) Value: %h\n", GRF6_26_buffer[clk]);
        end
        if (GRF6_27_buffer[clk] != GRF6_27_buffer[!clk]) begin
          $fwrite(f, "Register (6,27) Value: %h\n", GRF6_27_buffer[clk]);
        end
        if (GRF6_28_buffer[clk] != GRF6_28_buffer[!clk]) begin
          $fwrite(f, "Register (6,28) Value: %h\n", GRF6_28_buffer[clk]);
        end
        if (GRF6_29_buffer[clk] != GRF6_29_buffer[!clk]) begin
          $fwrite(f, "Register (6,29) Value: %h\n", GRF6_29_buffer[clk]);
        end
        if (GRF6_30_buffer[clk] != GRF6_30_buffer[!clk]) begin
          $fwrite(f, "Register (6,30) Value: %h\n", GRF6_30_buffer[clk]);
        end
        if (GRF6_31_buffer[clk] != GRF6_31_buffer[!clk]) begin
          $fwrite(f, "Register (6,31) Value: %h\n", GRF6_31_buffer[clk]);
        end
        if (GRF7_0_buffer[clk] != GRF7_0_buffer[!clk]) begin
          $fwrite(f, "Register (7,0) Value: %h\n", GRF7_0_buffer[clk]);
        end
        if (GRF7_1_buffer[clk] != GRF7_1_buffer[!clk]) begin
          $fwrite(f, "Register (7,1) Value: %h\n", GRF7_1_buffer[clk]);
        end
        if (GRF7_2_buffer[clk] != GRF7_2_buffer[!clk]) begin
          $fwrite(f, "Register (7,2) Value: %h\n", GRF7_2_buffer[clk]);
        end
        if (GRF7_3_buffer[clk] != GRF7_3_buffer[!clk]) begin
          $fwrite(f, "Register (7,3) Value: %h\n", GRF7_3_buffer[clk]);
        end
        if (GRF7_4_buffer[clk] != GRF7_4_buffer[!clk]) begin
          $fwrite(f, "Register (7,4) Value: %h\n", GRF7_4_buffer[clk]);
        end
        if (GRF7_5_buffer[clk] != GRF7_5_buffer[!clk]) begin
          $fwrite(f, "Register (7,5) Value: %h\n", GRF7_5_buffer[clk]);
        end
        if (GRF7_6_buffer[clk] != GRF7_6_buffer[!clk]) begin
          $fwrite(f, "Register (7,6) Value: %h\n", GRF7_6_buffer[clk]);
        end
        if (GRF7_7_buffer[clk] != GRF7_7_buffer[!clk]) begin
          $fwrite(f, "Register (7,7) Value: %h\n", GRF7_7_buffer[clk]);
        end
        if (GRF7_8_buffer[clk] != GRF7_8_buffer[!clk]) begin
          $fwrite(f, "Register (7,8) Value: %h\n", GRF7_8_buffer[clk]);
        end
        if (GRF7_9_buffer[clk] != GRF7_9_buffer[!clk]) begin
          $fwrite(f, "Register (7,9) Value: %h\n", GRF7_9_buffer[clk]);
        end
        if (GRF7_10_buffer[clk] != GRF7_10_buffer[!clk]) begin
          $fwrite(f, "Register (7,10) Value: %h\n", GRF7_10_buffer[clk]);
        end
        if (GRF7_11_buffer[clk] != GRF7_11_buffer[!clk]) begin
          $fwrite(f, "Register (7,11) Value: %h\n", GRF7_11_buffer[clk]);
        end
        if (GRF7_12_buffer[clk] != GRF7_12_buffer[!clk]) begin
          $fwrite(f, "Register (7,12) Value: %h\n", GRF7_12_buffer[clk]);
        end
        if (GRF7_13_buffer[clk] != GRF7_13_buffer[!clk]) begin
          $fwrite(f, "Register (7,13) Value: %h\n", GRF7_13_buffer[clk]);
        end
        if (GRF7_14_buffer[clk] != GRF7_14_buffer[!clk]) begin
          $fwrite(f, "Register (7,14) Value: %h\n", GRF7_14_buffer[clk]);
        end
        if (GRF7_15_buffer[clk] != GRF7_15_buffer[!clk]) begin
          $fwrite(f, "Register (7,15) Value: %h\n", GRF7_15_buffer[clk]);
        end
        if (GRF7_16_buffer[clk] != GRF7_16_buffer[!clk]) begin
          $fwrite(f, "Register (7,16) Value: %h\n", GRF7_16_buffer[clk]);
        end
        if (GRF7_17_buffer[clk] != GRF7_17_buffer[!clk]) begin
          $fwrite(f, "Register (7,17) Value: %h\n", GRF7_17_buffer[clk]);
        end
        if (GRF7_18_buffer[clk] != GRF7_18_buffer[!clk]) begin
          $fwrite(f, "Register (7,18) Value: %h\n", GRF7_18_buffer[clk]);
        end
        if (GRF7_19_buffer[clk] != GRF7_19_buffer[!clk]) begin
          $fwrite(f, "Register (7,19) Value: %h\n", GRF7_19_buffer[clk]);
        end
        if (GRF7_20_buffer[clk] != GRF7_20_buffer[!clk]) begin
          $fwrite(f, "Register (7,20) Value: %h\n", GRF7_20_buffer[clk]);
        end
        if (GRF7_21_buffer[clk] != GRF7_21_buffer[!clk]) begin
          $fwrite(f, "Register (7,21) Value: %h\n", GRF7_21_buffer[clk]);
        end
        if (GRF7_22_buffer[clk] != GRF7_22_buffer[!clk]) begin
          $fwrite(f, "Register (7,22) Value: %h\n", GRF7_22_buffer[clk]);
        end
        if (GRF7_23_buffer[clk] != GRF7_23_buffer[!clk]) begin
          $fwrite(f, "Register (7,23) Value: %h\n", GRF7_23_buffer[clk]);
        end
        if (GRF7_24_buffer[clk] != GRF7_24_buffer[!clk]) begin
          $fwrite(f, "Register (7,24) Value: %h\n", GRF7_24_buffer[clk]);
        end
        if (GRF7_25_buffer[clk] != GRF7_25_buffer[!clk]) begin
          $fwrite(f, "Register (7,25) Value: %h\n", GRF7_25_buffer[clk]);
        end
        if (GRF7_26_buffer[clk] != GRF7_26_buffer[!clk]) begin
          $fwrite(f, "Register (7,26) Value: %h\n", GRF7_26_buffer[clk]);
        end
        if (GRF7_27_buffer[clk] != GRF7_27_buffer[!clk]) begin
          $fwrite(f, "Register (7,27) Value: %h\n", GRF7_27_buffer[clk]);
        end
        if (GRF7_28_buffer[clk] != GRF7_28_buffer[!clk]) begin
          $fwrite(f, "Register (7,28) Value: %h\n", GRF7_28_buffer[clk]);
        end
        if (GRF7_29_buffer[clk] != GRF7_29_buffer[!clk]) begin
          $fwrite(f, "Register (7,29) Value: %h\n", GRF7_29_buffer[clk]);
        end
        if (GRF7_30_buffer[clk] != GRF7_30_buffer[!clk]) begin
          $fwrite(f, "Register (7,30) Value: %h\n", GRF7_30_buffer[clk]);
        end
        if (GRF7_31_buffer[clk] != GRF7_31_buffer[!clk]) begin
          $fwrite(f, "Register (7,31) Value: %h\n", GRF7_31_buffer[clk]);
        end
        if (GRF8_0_buffer[clk] != GRF8_0_buffer[!clk]) begin
          $fwrite(f, "Register (8,0) Value: %h\n", GRF8_0_buffer[clk]);
        end
        if (GRF8_1_buffer[clk] != GRF8_1_buffer[!clk]) begin
          $fwrite(f, "Register (8,1) Value: %h\n", GRF8_1_buffer[clk]);
        end
        if (GRF8_2_buffer[clk] != GRF8_2_buffer[!clk]) begin
          $fwrite(f, "Register (8,2) Value: %h\n", GRF8_2_buffer[clk]);
        end
        if (GRF8_3_buffer[clk] != GRF8_3_buffer[!clk]) begin
          $fwrite(f, "Register (8,3) Value: %h\n", GRF8_3_buffer[clk]);
        end
        if (GRF8_4_buffer[clk] != GRF8_4_buffer[!clk]) begin
          $fwrite(f, "Register (8,4) Value: %h\n", GRF8_4_buffer[clk]);
        end
        if (GRF8_5_buffer[clk] != GRF8_5_buffer[!clk]) begin
          $fwrite(f, "Register (8,5) Value: %h\n", GRF8_5_buffer[clk]);
        end
        if (GRF8_6_buffer[clk] != GRF8_6_buffer[!clk]) begin
          $fwrite(f, "Register (8,6) Value: %h\n", GRF8_6_buffer[clk]);
        end
        if (GRF8_7_buffer[clk] != GRF8_7_buffer[!clk]) begin
          $fwrite(f, "Register (8,7) Value: %h\n", GRF8_7_buffer[clk]);
        end
        if (GRF8_8_buffer[clk] != GRF8_8_buffer[!clk]) begin
          $fwrite(f, "Register (8,8) Value: %h\n", GRF8_8_buffer[clk]);
        end
        if (GRF8_9_buffer[clk] != GRF8_9_buffer[!clk]) begin
          $fwrite(f, "Register (8,9) Value: %h\n", GRF8_9_buffer[clk]);
        end
        if (GRF8_10_buffer[clk] != GRF8_10_buffer[!clk]) begin
          $fwrite(f, "Register (8,10) Value: %h\n", GRF8_10_buffer[clk]);
        end
        if (GRF8_11_buffer[clk] != GRF8_11_buffer[!clk]) begin
          $fwrite(f, "Register (8,11) Value: %h\n", GRF8_11_buffer[clk]);
        end
        if (GRF8_12_buffer[clk] != GRF8_12_buffer[!clk]) begin
          $fwrite(f, "Register (8,12) Value: %h\n", GRF8_12_buffer[clk]);
        end
        if (GRF8_13_buffer[clk] != GRF8_13_buffer[!clk]) begin
          $fwrite(f, "Register (8,13) Value: %h\n", GRF8_13_buffer[clk]);
        end
        if (GRF8_14_buffer[clk] != GRF8_14_buffer[!clk]) begin
          $fwrite(f, "Register (8,14) Value: %h\n", GRF8_14_buffer[clk]);
        end
        if (GRF8_15_buffer[clk] != GRF8_15_buffer[!clk]) begin
          $fwrite(f, "Register (8,15) Value: %h\n", GRF8_15_buffer[clk]);
        end
        if (GRF8_16_buffer[clk] != GRF8_16_buffer[!clk]) begin
          $fwrite(f, "Register (8,16) Value: %h\n", GRF8_16_buffer[clk]);
        end
        if (GRF8_17_buffer[clk] != GRF8_17_buffer[!clk]) begin
          $fwrite(f, "Register (8,17) Value: %h\n", GRF8_17_buffer[clk]);
        end
        if (GRF8_18_buffer[clk] != GRF8_18_buffer[!clk]) begin
          $fwrite(f, "Register (8,18) Value: %h\n", GRF8_18_buffer[clk]);
        end
        if (GRF8_19_buffer[clk] != GRF8_19_buffer[!clk]) begin
          $fwrite(f, "Register (8,19) Value: %h\n", GRF8_19_buffer[clk]);
        end
        if (GRF8_20_buffer[clk] != GRF8_20_buffer[!clk]) begin
          $fwrite(f, "Register (8,20) Value: %h\n", GRF8_20_buffer[clk]);
        end
        if (GRF8_21_buffer[clk] != GRF8_21_buffer[!clk]) begin
          $fwrite(f, "Register (8,21) Value: %h\n", GRF8_21_buffer[clk]);
        end
        if (GRF8_22_buffer[clk] != GRF8_22_buffer[!clk]) begin
          $fwrite(f, "Register (8,22) Value: %h\n", GRF8_22_buffer[clk]);
        end
        if (GRF8_23_buffer[clk] != GRF8_23_buffer[!clk]) begin
          $fwrite(f, "Register (8,23) Value: %h\n", GRF8_23_buffer[clk]);
        end
        if (GRF8_24_buffer[clk] != GRF8_24_buffer[!clk]) begin
          $fwrite(f, "Register (8,24) Value: %h\n", GRF8_24_buffer[clk]);
        end
        if (GRF8_25_buffer[clk] != GRF8_25_buffer[!clk]) begin
          $fwrite(f, "Register (8,25) Value: %h\n", GRF8_25_buffer[clk]);
        end
        if (GRF8_26_buffer[clk] != GRF8_26_buffer[!clk]) begin
          $fwrite(f, "Register (8,26) Value: %h\n", GRF8_26_buffer[clk]);
        end
        if (GRF8_27_buffer[clk] != GRF8_27_buffer[!clk]) begin
          $fwrite(f, "Register (8,27) Value: %h\n", GRF8_27_buffer[clk]);
        end
        if (GRF8_28_buffer[clk] != GRF8_28_buffer[!clk]) begin
          $fwrite(f, "Register (8,28) Value: %h\n", GRF8_28_buffer[clk]);
        end
        if (GRF8_29_buffer[clk] != GRF8_29_buffer[!clk]) begin
          $fwrite(f, "Register (8,29) Value: %h\n", GRF8_29_buffer[clk]);
        end
        if (GRF8_30_buffer[clk] != GRF8_30_buffer[!clk]) begin
          $fwrite(f, "Register (8,30) Value: %h\n", GRF8_30_buffer[clk]);
        end
        if (GRF8_31_buffer[clk] != GRF8_31_buffer[!clk]) begin
          $fwrite(f, "Register (8,31) Value: %h\n", GRF8_31_buffer[clk]);
        end
        if (GRF9_0_buffer[clk] != GRF9_0_buffer[!clk]) begin
          $fwrite(f, "Register (9,0) Value: %h\n", GRF9_0_buffer[clk]);
        end
        if (GRF9_1_buffer[clk] != GRF9_1_buffer[!clk]) begin
          $fwrite(f, "Register (9,1) Value: %h\n", GRF9_1_buffer[clk]);
        end
        if (GRF9_2_buffer[clk] != GRF9_2_buffer[!clk]) begin
          $fwrite(f, "Register (9,2) Value: %h\n", GRF9_2_buffer[clk]);
        end
        if (GRF9_3_buffer[clk] != GRF9_3_buffer[!clk]) begin
          $fwrite(f, "Register (9,3) Value: %h\n", GRF9_3_buffer[clk]);
        end
        if (GRF9_4_buffer[clk] != GRF9_4_buffer[!clk]) begin
          $fwrite(f, "Register (9,4) Value: %h\n", GRF9_4_buffer[clk]);
        end
        if (GRF9_5_buffer[clk] != GRF9_5_buffer[!clk]) begin
          $fwrite(f, "Register (9,5) Value: %h\n", GRF9_5_buffer[clk]);
        end
        if (GRF9_6_buffer[clk] != GRF9_6_buffer[!clk]) begin
          $fwrite(f, "Register (9,6) Value: %h\n", GRF9_6_buffer[clk]);
        end
        if (GRF9_7_buffer[clk] != GRF9_7_buffer[!clk]) begin
          $fwrite(f, "Register (9,7) Value: %h\n", GRF9_7_buffer[clk]);
        end
        if (GRF9_8_buffer[clk] != GRF9_8_buffer[!clk]) begin
          $fwrite(f, "Register (9,8) Value: %h\n", GRF9_8_buffer[clk]);
        end
        if (GRF9_9_buffer[clk] != GRF9_9_buffer[!clk]) begin
          $fwrite(f, "Register (9,9) Value: %h\n", GRF9_9_buffer[clk]);
        end
        if (GRF9_10_buffer[clk] != GRF9_10_buffer[!clk]) begin
          $fwrite(f, "Register (9,10) Value: %h\n", GRF9_10_buffer[clk]);
        end
        if (GRF9_11_buffer[clk] != GRF9_11_buffer[!clk]) begin
          $fwrite(f, "Register (9,11) Value: %h\n", GRF9_11_buffer[clk]);
        end
        if (GRF9_12_buffer[clk] != GRF9_12_buffer[!clk]) begin
          $fwrite(f, "Register (9,12) Value: %h\n", GRF9_12_buffer[clk]);
        end
        if (GRF9_13_buffer[clk] != GRF9_13_buffer[!clk]) begin
          $fwrite(f, "Register (9,13) Value: %h\n", GRF9_13_buffer[clk]);
        end
        if (GRF9_14_buffer[clk] != GRF9_14_buffer[!clk]) begin
          $fwrite(f, "Register (9,14) Value: %h\n", GRF9_14_buffer[clk]);
        end
        if (GRF9_15_buffer[clk] != GRF9_15_buffer[!clk]) begin
          $fwrite(f, "Register (9,15) Value: %h\n", GRF9_15_buffer[clk]);
        end
        if (GRF9_16_buffer[clk] != GRF9_16_buffer[!clk]) begin
          $fwrite(f, "Register (9,16) Value: %h\n", GRF9_16_buffer[clk]);
        end
        if (GRF9_17_buffer[clk] != GRF9_17_buffer[!clk]) begin
          $fwrite(f, "Register (9,17) Value: %h\n", GRF9_17_buffer[clk]);
        end
        if (GRF9_18_buffer[clk] != GRF9_18_buffer[!clk]) begin
          $fwrite(f, "Register (9,18) Value: %h\n", GRF9_18_buffer[clk]);
        end
        if (GRF9_19_buffer[clk] != GRF9_19_buffer[!clk]) begin
          $fwrite(f, "Register (9,19) Value: %h\n", GRF9_19_buffer[clk]);
        end
        if (GRF9_20_buffer[clk] != GRF9_20_buffer[!clk]) begin
          $fwrite(f, "Register (9,20) Value: %h\n", GRF9_20_buffer[clk]);
        end
        if (GRF9_21_buffer[clk] != GRF9_21_buffer[!clk]) begin
          $fwrite(f, "Register (9,21) Value: %h\n", GRF9_21_buffer[clk]);
        end
        if (GRF9_22_buffer[clk] != GRF9_22_buffer[!clk]) begin
          $fwrite(f, "Register (9,22) Value: %h\n", GRF9_22_buffer[clk]);
        end
        if (GRF9_23_buffer[clk] != GRF9_23_buffer[!clk]) begin
          $fwrite(f, "Register (9,23) Value: %h\n", GRF9_23_buffer[clk]);
        end
        if (GRF9_24_buffer[clk] != GRF9_24_buffer[!clk]) begin
          $fwrite(f, "Register (9,24) Value: %h\n", GRF9_24_buffer[clk]);
        end
        if (GRF9_25_buffer[clk] != GRF9_25_buffer[!clk]) begin
          $fwrite(f, "Register (9,25) Value: %h\n", GRF9_25_buffer[clk]);
        end
        if (GRF9_26_buffer[clk] != GRF9_26_buffer[!clk]) begin
          $fwrite(f, "Register (9,26) Value: %h\n", GRF9_26_buffer[clk]);
        end
        if (GRF9_27_buffer[clk] != GRF9_27_buffer[!clk]) begin
          $fwrite(f, "Register (9,27) Value: %h\n", GRF9_27_buffer[clk]);
        end
        if (GRF9_28_buffer[clk] != GRF9_28_buffer[!clk]) begin
          $fwrite(f, "Register (9,28) Value: %h\n", GRF9_28_buffer[clk]);
        end
        if (GRF9_29_buffer[clk] != GRF9_29_buffer[!clk]) begin
          $fwrite(f, "Register (9,29) Value: %h\n", GRF9_29_buffer[clk]);
        end
        if (GRF9_30_buffer[clk] != GRF9_30_buffer[!clk]) begin
          $fwrite(f, "Register (9,30) Value: %h\n", GRF9_30_buffer[clk]);
        end
        if (GRF9_31_buffer[clk] != GRF9_31_buffer[!clk]) begin
          $fwrite(f, "Register (9,31) Value: %h\n", GRF9_31_buffer[clk]);
        end
        if (GRF10_0_buffer[clk] != GRF10_0_buffer[!clk]) begin
          $fwrite(f, "Register (10,0) Value: %h\n", GRF10_0_buffer[clk]);
        end
        if (GRF10_1_buffer[clk] != GRF10_1_buffer[!clk]) begin
          $fwrite(f, "Register (10,1) Value: %h\n", GRF10_1_buffer[clk]);
        end
        if (GRF10_2_buffer[clk] != GRF10_2_buffer[!clk]) begin
          $fwrite(f, "Register (10,2) Value: %h\n", GRF10_2_buffer[clk]);
        end
        if (GRF10_3_buffer[clk] != GRF10_3_buffer[!clk]) begin
          $fwrite(f, "Register (10,3) Value: %h\n", GRF10_3_buffer[clk]);
        end
        if (GRF10_4_buffer[clk] != GRF10_4_buffer[!clk]) begin
          $fwrite(f, "Register (10,4) Value: %h\n", GRF10_4_buffer[clk]);
        end
        if (GRF10_5_buffer[clk] != GRF10_5_buffer[!clk]) begin
          $fwrite(f, "Register (10,5) Value: %h\n", GRF10_5_buffer[clk]);
        end
        if (GRF10_6_buffer[clk] != GRF10_6_buffer[!clk]) begin
          $fwrite(f, "Register (10,6) Value: %h\n", GRF10_6_buffer[clk]);
        end
        if (GRF10_7_buffer[clk] != GRF10_7_buffer[!clk]) begin
          $fwrite(f, "Register (10,7) Value: %h\n", GRF10_7_buffer[clk]);
        end
        if (GRF10_8_buffer[clk] != GRF10_8_buffer[!clk]) begin
          $fwrite(f, "Register (10,8) Value: %h\n", GRF10_8_buffer[clk]);
        end
        if (GRF10_9_buffer[clk] != GRF10_9_buffer[!clk]) begin
          $fwrite(f, "Register (10,9) Value: %h\n", GRF10_9_buffer[clk]);
        end
        if (GRF10_10_buffer[clk] != GRF10_10_buffer[!clk]) begin
          $fwrite(f, "Register (10,10) Value: %h\n", GRF10_10_buffer[clk]);
        end
        if (GRF10_11_buffer[clk] != GRF10_11_buffer[!clk]) begin
          $fwrite(f, "Register (10,11) Value: %h\n", GRF10_11_buffer[clk]);
        end
        if (GRF10_12_buffer[clk] != GRF10_12_buffer[!clk]) begin
          $fwrite(f, "Register (10,12) Value: %h\n", GRF10_12_buffer[clk]);
        end
        if (GRF10_13_buffer[clk] != GRF10_13_buffer[!clk]) begin
          $fwrite(f, "Register (10,13) Value: %h\n", GRF10_13_buffer[clk]);
        end
        if (GRF10_14_buffer[clk] != GRF10_14_buffer[!clk]) begin
          $fwrite(f, "Register (10,14) Value: %h\n", GRF10_14_buffer[clk]);
        end
        if (GRF10_15_buffer[clk] != GRF10_15_buffer[!clk]) begin
          $fwrite(f, "Register (10,15) Value: %h\n", GRF10_15_buffer[clk]);
        end
        if (GRF10_16_buffer[clk] != GRF10_16_buffer[!clk]) begin
          $fwrite(f, "Register (10,16) Value: %h\n", GRF10_16_buffer[clk]);
        end
        if (GRF10_17_buffer[clk] != GRF10_17_buffer[!clk]) begin
          $fwrite(f, "Register (10,17) Value: %h\n", GRF10_17_buffer[clk]);
        end
        if (GRF10_18_buffer[clk] != GRF10_18_buffer[!clk]) begin
          $fwrite(f, "Register (10,18) Value: %h\n", GRF10_18_buffer[clk]);
        end
        if (GRF10_19_buffer[clk] != GRF10_19_buffer[!clk]) begin
          $fwrite(f, "Register (10,19) Value: %h\n", GRF10_19_buffer[clk]);
        end
        if (GRF10_20_buffer[clk] != GRF10_20_buffer[!clk]) begin
          $fwrite(f, "Register (10,20) Value: %h\n", GRF10_20_buffer[clk]);
        end
        if (GRF10_21_buffer[clk] != GRF10_21_buffer[!clk]) begin
          $fwrite(f, "Register (10,21) Value: %h\n", GRF10_21_buffer[clk]);
        end
        if (GRF10_22_buffer[clk] != GRF10_22_buffer[!clk]) begin
          $fwrite(f, "Register (10,22) Value: %h\n", GRF10_22_buffer[clk]);
        end
        if (GRF10_23_buffer[clk] != GRF10_23_buffer[!clk]) begin
          $fwrite(f, "Register (10,23) Value: %h\n", GRF10_23_buffer[clk]);
        end
        if (GRF10_24_buffer[clk] != GRF10_24_buffer[!clk]) begin
          $fwrite(f, "Register (10,24) Value: %h\n", GRF10_24_buffer[clk]);
        end
        if (GRF10_25_buffer[clk] != GRF10_25_buffer[!clk]) begin
          $fwrite(f, "Register (10,25) Value: %h\n", GRF10_25_buffer[clk]);
        end
        if (GRF10_26_buffer[clk] != GRF10_26_buffer[!clk]) begin
          $fwrite(f, "Register (10,26) Value: %h\n", GRF10_26_buffer[clk]);
        end
        if (GRF10_27_buffer[clk] != GRF10_27_buffer[!clk]) begin
          $fwrite(f, "Register (10,27) Value: %h\n", GRF10_27_buffer[clk]);
        end
        if (GRF10_28_buffer[clk] != GRF10_28_buffer[!clk]) begin
          $fwrite(f, "Register (10,28) Value: %h\n", GRF10_28_buffer[clk]);
        end
        if (GRF10_29_buffer[clk] != GRF10_29_buffer[!clk]) begin
          $fwrite(f, "Register (10,29) Value: %h\n", GRF10_29_buffer[clk]);
        end
        if (GRF10_30_buffer[clk] != GRF10_30_buffer[!clk]) begin
          $fwrite(f, "Register (10,30) Value: %h\n", GRF10_30_buffer[clk]);
        end
        if (GRF10_31_buffer[clk] != GRF10_31_buffer[!clk]) begin
          $fwrite(f, "Register (10,31) Value: %h\n", GRF10_31_buffer[clk]);
        end
        if (GRF11_0_buffer[clk] != GRF11_0_buffer[!clk]) begin
          $fwrite(f, "Register (11,0) Value: %h\n", GRF11_0_buffer[clk]);
        end
        if (GRF11_1_buffer[clk] != GRF11_1_buffer[!clk]) begin
          $fwrite(f, "Register (11,1) Value: %h\n", GRF11_1_buffer[clk]);
        end
        if (GRF11_2_buffer[clk] != GRF11_2_buffer[!clk]) begin
          $fwrite(f, "Register (11,2) Value: %h\n", GRF11_2_buffer[clk]);
        end
        if (GRF11_3_buffer[clk] != GRF11_3_buffer[!clk]) begin
          $fwrite(f, "Register (11,3) Value: %h\n", GRF11_3_buffer[clk]);
        end
        if (GRF11_4_buffer[clk] != GRF11_4_buffer[!clk]) begin
          $fwrite(f, "Register (11,4) Value: %h\n", GRF11_4_buffer[clk]);
        end
        if (GRF11_5_buffer[clk] != GRF11_5_buffer[!clk]) begin
          $fwrite(f, "Register (11,5) Value: %h\n", GRF11_5_buffer[clk]);
        end
        if (GRF11_6_buffer[clk] != GRF11_6_buffer[!clk]) begin
          $fwrite(f, "Register (11,6) Value: %h\n", GRF11_6_buffer[clk]);
        end
        if (GRF11_7_buffer[clk] != GRF11_7_buffer[!clk]) begin
          $fwrite(f, "Register (11,7) Value: %h\n", GRF11_7_buffer[clk]);
        end
        if (GRF11_8_buffer[clk] != GRF11_8_buffer[!clk]) begin
          $fwrite(f, "Register (11,8) Value: %h\n", GRF11_8_buffer[clk]);
        end
        if (GRF11_9_buffer[clk] != GRF11_9_buffer[!clk]) begin
          $fwrite(f, "Register (11,9) Value: %h\n", GRF11_9_buffer[clk]);
        end
        if (GRF11_10_buffer[clk] != GRF11_10_buffer[!clk]) begin
          $fwrite(f, "Register (11,10) Value: %h\n", GRF11_10_buffer[clk]);
        end
        if (GRF11_11_buffer[clk] != GRF11_11_buffer[!clk]) begin
          $fwrite(f, "Register (11,11) Value: %h\n", GRF11_11_buffer[clk]);
        end
        if (GRF11_12_buffer[clk] != GRF11_12_buffer[!clk]) begin
          $fwrite(f, "Register (11,12) Value: %h\n", GRF11_12_buffer[clk]);
        end
        if (GRF11_13_buffer[clk] != GRF11_13_buffer[!clk]) begin
          $fwrite(f, "Register (11,13) Value: %h\n", GRF11_13_buffer[clk]);
        end
        if (GRF11_14_buffer[clk] != GRF11_14_buffer[!clk]) begin
          $fwrite(f, "Register (11,14) Value: %h\n", GRF11_14_buffer[clk]);
        end
        if (GRF11_15_buffer[clk] != GRF11_15_buffer[!clk]) begin
          $fwrite(f, "Register (11,15) Value: %h\n", GRF11_15_buffer[clk]);
        end
        if (GRF11_16_buffer[clk] != GRF11_16_buffer[!clk]) begin
          $fwrite(f, "Register (11,16) Value: %h\n", GRF11_16_buffer[clk]);
        end
        if (GRF11_17_buffer[clk] != GRF11_17_buffer[!clk]) begin
          $fwrite(f, "Register (11,17) Value: %h\n", GRF11_17_buffer[clk]);
        end
        if (GRF11_18_buffer[clk] != GRF11_18_buffer[!clk]) begin
          $fwrite(f, "Register (11,18) Value: %h\n", GRF11_18_buffer[clk]);
        end
        if (GRF11_19_buffer[clk] != GRF11_19_buffer[!clk]) begin
          $fwrite(f, "Register (11,19) Value: %h\n", GRF11_19_buffer[clk]);
        end
        if (GRF11_20_buffer[clk] != GRF11_20_buffer[!clk]) begin
          $fwrite(f, "Register (11,20) Value: %h\n", GRF11_20_buffer[clk]);
        end
        if (GRF11_21_buffer[clk] != GRF11_21_buffer[!clk]) begin
          $fwrite(f, "Register (11,21) Value: %h\n", GRF11_21_buffer[clk]);
        end
        if (GRF11_22_buffer[clk] != GRF11_22_buffer[!clk]) begin
          $fwrite(f, "Register (11,22) Value: %h\n", GRF11_22_buffer[clk]);
        end
        if (GRF11_23_buffer[clk] != GRF11_23_buffer[!clk]) begin
          $fwrite(f, "Register (11,23) Value: %h\n", GRF11_23_buffer[clk]);
        end
        if (GRF11_24_buffer[clk] != GRF11_24_buffer[!clk]) begin
          $fwrite(f, "Register (11,24) Value: %h\n", GRF11_24_buffer[clk]);
        end
        if (GRF11_25_buffer[clk] != GRF11_25_buffer[!clk]) begin
          $fwrite(f, "Register (11,25) Value: %h\n", GRF11_25_buffer[clk]);
        end
        if (GRF11_26_buffer[clk] != GRF11_26_buffer[!clk]) begin
          $fwrite(f, "Register (11,26) Value: %h\n", GRF11_26_buffer[clk]);
        end
        if (GRF11_27_buffer[clk] != GRF11_27_buffer[!clk]) begin
          $fwrite(f, "Register (11,27) Value: %h\n", GRF11_27_buffer[clk]);
        end
        if (GRF11_28_buffer[clk] != GRF11_28_buffer[!clk]) begin
          $fwrite(f, "Register (11,28) Value: %h\n", GRF11_28_buffer[clk]);
        end
        if (GRF11_29_buffer[clk] != GRF11_29_buffer[!clk]) begin
          $fwrite(f, "Register (11,29) Value: %h\n", GRF11_29_buffer[clk]);
        end
        if (GRF11_30_buffer[clk] != GRF11_30_buffer[!clk]) begin
          $fwrite(f, "Register (11,30) Value: %h\n", GRF11_30_buffer[clk]);
        end
        if (GRF11_31_buffer[clk] != GRF11_31_buffer[!clk]) begin
          $fwrite(f, "Register (11,31) Value: %h\n", GRF11_31_buffer[clk]);
        end
        if (GRF12_0_buffer[clk] != GRF12_0_buffer[!clk]) begin
          $fwrite(f, "Register (12,0) Value: %h\n", GRF12_0_buffer[clk]);
        end
        if (GRF12_1_buffer[clk] != GRF12_1_buffer[!clk]) begin
          $fwrite(f, "Register (12,1) Value: %h\n", GRF12_1_buffer[clk]);
        end
        if (GRF12_2_buffer[clk] != GRF12_2_buffer[!clk]) begin
          $fwrite(f, "Register (12,2) Value: %h\n", GRF12_2_buffer[clk]);
        end
        if (GRF12_3_buffer[clk] != GRF12_3_buffer[!clk]) begin
          $fwrite(f, "Register (12,3) Value: %h\n", GRF12_3_buffer[clk]);
        end
        if (GRF12_4_buffer[clk] != GRF12_4_buffer[!clk]) begin
          $fwrite(f, "Register (12,4) Value: %h\n", GRF12_4_buffer[clk]);
        end
        if (GRF12_5_buffer[clk] != GRF12_5_buffer[!clk]) begin
          $fwrite(f, "Register (12,5) Value: %h\n", GRF12_5_buffer[clk]);
        end
        if (GRF12_6_buffer[clk] != GRF12_6_buffer[!clk]) begin
          $fwrite(f, "Register (12,6) Value: %h\n", GRF12_6_buffer[clk]);
        end
        if (GRF12_7_buffer[clk] != GRF12_7_buffer[!clk]) begin
          $fwrite(f, "Register (12,7) Value: %h\n", GRF12_7_buffer[clk]);
        end
        if (GRF12_8_buffer[clk] != GRF12_8_buffer[!clk]) begin
          $fwrite(f, "Register (12,8) Value: %h\n", GRF12_8_buffer[clk]);
        end
        if (GRF12_9_buffer[clk] != GRF12_9_buffer[!clk]) begin
          $fwrite(f, "Register (12,9) Value: %h\n", GRF12_9_buffer[clk]);
        end
        if (GRF12_10_buffer[clk] != GRF12_10_buffer[!clk]) begin
          $fwrite(f, "Register (12,10) Value: %h\n", GRF12_10_buffer[clk]);
        end
        if (GRF12_11_buffer[clk] != GRF12_11_buffer[!clk]) begin
          $fwrite(f, "Register (12,11) Value: %h\n", GRF12_11_buffer[clk]);
        end
        if (GRF12_12_buffer[clk] != GRF12_12_buffer[!clk]) begin
          $fwrite(f, "Register (12,12) Value: %h\n", GRF12_12_buffer[clk]);
        end
        if (GRF12_13_buffer[clk] != GRF12_13_buffer[!clk]) begin
          $fwrite(f, "Register (12,13) Value: %h\n", GRF12_13_buffer[clk]);
        end
        if (GRF12_14_buffer[clk] != GRF12_14_buffer[!clk]) begin
          $fwrite(f, "Register (12,14) Value: %h\n", GRF12_14_buffer[clk]);
        end
        if (GRF12_15_buffer[clk] != GRF12_15_buffer[!clk]) begin
          $fwrite(f, "Register (12,15) Value: %h\n", GRF12_15_buffer[clk]);
        end
        if (GRF12_16_buffer[clk] != GRF12_16_buffer[!clk]) begin
          $fwrite(f, "Register (12,16) Value: %h\n", GRF12_16_buffer[clk]);
        end
        if (GRF12_17_buffer[clk] != GRF12_17_buffer[!clk]) begin
          $fwrite(f, "Register (12,17) Value: %h\n", GRF12_17_buffer[clk]);
        end
        if (GRF12_18_buffer[clk] != GRF12_18_buffer[!clk]) begin
          $fwrite(f, "Register (12,18) Value: %h\n", GRF12_18_buffer[clk]);
        end
        if (GRF12_19_buffer[clk] != GRF12_19_buffer[!clk]) begin
          $fwrite(f, "Register (12,19) Value: %h\n", GRF12_19_buffer[clk]);
        end
        if (GRF12_20_buffer[clk] != GRF12_20_buffer[!clk]) begin
          $fwrite(f, "Register (12,20) Value: %h\n", GRF12_20_buffer[clk]);
        end
        if (GRF12_21_buffer[clk] != GRF12_21_buffer[!clk]) begin
          $fwrite(f, "Register (12,21) Value: %h\n", GRF12_21_buffer[clk]);
        end
        if (GRF12_22_buffer[clk] != GRF12_22_buffer[!clk]) begin
          $fwrite(f, "Register (12,22) Value: %h\n", GRF12_22_buffer[clk]);
        end
        if (GRF12_23_buffer[clk] != GRF12_23_buffer[!clk]) begin
          $fwrite(f, "Register (12,23) Value: %h\n", GRF12_23_buffer[clk]);
        end
        if (GRF12_24_buffer[clk] != GRF12_24_buffer[!clk]) begin
          $fwrite(f, "Register (12,24) Value: %h\n", GRF12_24_buffer[clk]);
        end
        if (GRF12_25_buffer[clk] != GRF12_25_buffer[!clk]) begin
          $fwrite(f, "Register (12,25) Value: %h\n", GRF12_25_buffer[clk]);
        end
        if (GRF12_26_buffer[clk] != GRF12_26_buffer[!clk]) begin
          $fwrite(f, "Register (12,26) Value: %h\n", GRF12_26_buffer[clk]);
        end
        if (GRF12_27_buffer[clk] != GRF12_27_buffer[!clk]) begin
          $fwrite(f, "Register (12,27) Value: %h\n", GRF12_27_buffer[clk]);
        end
        if (GRF12_28_buffer[clk] != GRF12_28_buffer[!clk]) begin
          $fwrite(f, "Register (12,28) Value: %h\n", GRF12_28_buffer[clk]);
        end
        if (GRF12_29_buffer[clk] != GRF12_29_buffer[!clk]) begin
          $fwrite(f, "Register (12,29) Value: %h\n", GRF12_29_buffer[clk]);
        end
        if (GRF12_30_buffer[clk] != GRF12_30_buffer[!clk]) begin
          $fwrite(f, "Register (12,30) Value: %h\n", GRF12_30_buffer[clk]);
        end
        if (GRF12_31_buffer[clk] != GRF12_31_buffer[!clk]) begin
          $fwrite(f, "Register (12,31) Value: %h\n", GRF12_31_buffer[clk]);
        end
        if (GRF13_0_buffer[clk] != GRF13_0_buffer[!clk]) begin
          $fwrite(f, "Register (13,0) Value: %h\n", GRF13_0_buffer[clk]);
        end
        if (GRF13_1_buffer[clk] != GRF13_1_buffer[!clk]) begin
          $fwrite(f, "Register (13,1) Value: %h\n", GRF13_1_buffer[clk]);
        end
        if (GRF13_2_buffer[clk] != GRF13_2_buffer[!clk]) begin
          $fwrite(f, "Register (13,2) Value: %h\n", GRF13_2_buffer[clk]);
        end
        if (GRF13_3_buffer[clk] != GRF13_3_buffer[!clk]) begin
          $fwrite(f, "Register (13,3) Value: %h\n", GRF13_3_buffer[clk]);
        end
        if (GRF13_4_buffer[clk] != GRF13_4_buffer[!clk]) begin
          $fwrite(f, "Register (13,4) Value: %h\n", GRF13_4_buffer[clk]);
        end
        if (GRF13_5_buffer[clk] != GRF13_5_buffer[!clk]) begin
          $fwrite(f, "Register (13,5) Value: %h\n", GRF13_5_buffer[clk]);
        end
        if (GRF13_6_buffer[clk] != GRF13_6_buffer[!clk]) begin
          $fwrite(f, "Register (13,6) Value: %h\n", GRF13_6_buffer[clk]);
        end
        if (GRF13_7_buffer[clk] != GRF13_7_buffer[!clk]) begin
          $fwrite(f, "Register (13,7) Value: %h\n", GRF13_7_buffer[clk]);
        end
        if (GRF13_8_buffer[clk] != GRF13_8_buffer[!clk]) begin
          $fwrite(f, "Register (13,8) Value: %h\n", GRF13_8_buffer[clk]);
        end
        if (GRF13_9_buffer[clk] != GRF13_9_buffer[!clk]) begin
          $fwrite(f, "Register (13,9) Value: %h\n", GRF13_9_buffer[clk]);
        end
        if (GRF13_10_buffer[clk] != GRF13_10_buffer[!clk]) begin
          $fwrite(f, "Register (13,10) Value: %h\n", GRF13_10_buffer[clk]);
        end
        if (GRF13_11_buffer[clk] != GRF13_11_buffer[!clk]) begin
          $fwrite(f, "Register (13,11) Value: %h\n", GRF13_11_buffer[clk]);
        end
        if (GRF13_12_buffer[clk] != GRF13_12_buffer[!clk]) begin
          $fwrite(f, "Register (13,12) Value: %h\n", GRF13_12_buffer[clk]);
        end
        if (GRF13_13_buffer[clk] != GRF13_13_buffer[!clk]) begin
          $fwrite(f, "Register (13,13) Value: %h\n", GRF13_13_buffer[clk]);
        end
        if (GRF13_14_buffer[clk] != GRF13_14_buffer[!clk]) begin
          $fwrite(f, "Register (13,14) Value: %h\n", GRF13_14_buffer[clk]);
        end
        if (GRF13_15_buffer[clk] != GRF13_15_buffer[!clk]) begin
          $fwrite(f, "Register (13,15) Value: %h\n", GRF13_15_buffer[clk]);
        end
        if (GRF13_16_buffer[clk] != GRF13_16_buffer[!clk]) begin
          $fwrite(f, "Register (13,16) Value: %h\n", GRF13_16_buffer[clk]);
        end
        if (GRF13_17_buffer[clk] != GRF13_17_buffer[!clk]) begin
          $fwrite(f, "Register (13,17) Value: %h\n", GRF13_17_buffer[clk]);
        end
        if (GRF13_18_buffer[clk] != GRF13_18_buffer[!clk]) begin
          $fwrite(f, "Register (13,18) Value: %h\n", GRF13_18_buffer[clk]);
        end
        if (GRF13_19_buffer[clk] != GRF13_19_buffer[!clk]) begin
          $fwrite(f, "Register (13,19) Value: %h\n", GRF13_19_buffer[clk]);
        end
        if (GRF13_20_buffer[clk] != GRF13_20_buffer[!clk]) begin
          $fwrite(f, "Register (13,20) Value: %h\n", GRF13_20_buffer[clk]);
        end
        if (GRF13_21_buffer[clk] != GRF13_21_buffer[!clk]) begin
          $fwrite(f, "Register (13,21) Value: %h\n", GRF13_21_buffer[clk]);
        end
        if (GRF13_22_buffer[clk] != GRF13_22_buffer[!clk]) begin
          $fwrite(f, "Register (13,22) Value: %h\n", GRF13_22_buffer[clk]);
        end
        if (GRF13_23_buffer[clk] != GRF13_23_buffer[!clk]) begin
          $fwrite(f, "Register (13,23) Value: %h\n", GRF13_23_buffer[clk]);
        end
        if (GRF13_24_buffer[clk] != GRF13_24_buffer[!clk]) begin
          $fwrite(f, "Register (13,24) Value: %h\n", GRF13_24_buffer[clk]);
        end
        if (GRF13_25_buffer[clk] != GRF13_25_buffer[!clk]) begin
          $fwrite(f, "Register (13,25) Value: %h\n", GRF13_25_buffer[clk]);
        end
        if (GRF13_26_buffer[clk] != GRF13_26_buffer[!clk]) begin
          $fwrite(f, "Register (13,26) Value: %h\n", GRF13_26_buffer[clk]);
        end
        if (GRF13_27_buffer[clk] != GRF13_27_buffer[!clk]) begin
          $fwrite(f, "Register (13,27) Value: %h\n", GRF13_27_buffer[clk]);
        end
        if (GRF13_28_buffer[clk] != GRF13_28_buffer[!clk]) begin
          $fwrite(f, "Register (13,28) Value: %h\n", GRF13_28_buffer[clk]);
        end
        if (GRF13_29_buffer[clk] != GRF13_29_buffer[!clk]) begin
          $fwrite(f, "Register (13,29) Value: %h\n", GRF13_29_buffer[clk]);
        end
        if (GRF13_30_buffer[clk] != GRF13_30_buffer[!clk]) begin
          $fwrite(f, "Register (13,30) Value: %h\n", GRF13_30_buffer[clk]);
        end
        if (GRF13_31_buffer[clk] != GRF13_31_buffer[!clk]) begin
          $fwrite(f, "Register (13,31) Value: %h\n", GRF13_31_buffer[clk]);
        end
        if (GRF14_0_buffer[clk] != GRF14_0_buffer[!clk]) begin
          $fwrite(f, "Register (14,0) Value: %h\n", GRF14_0_buffer[clk]);
        end
        if (GRF14_1_buffer[clk] != GRF14_1_buffer[!clk]) begin
          $fwrite(f, "Register (14,1) Value: %h\n", GRF14_1_buffer[clk]);
        end
        if (GRF14_2_buffer[clk] != GRF14_2_buffer[!clk]) begin
          $fwrite(f, "Register (14,2) Value: %h\n", GRF14_2_buffer[clk]);
        end
        if (GRF14_3_buffer[clk] != GRF14_3_buffer[!clk]) begin
          $fwrite(f, "Register (14,3) Value: %h\n", GRF14_3_buffer[clk]);
        end
        if (GRF14_4_buffer[clk] != GRF14_4_buffer[!clk]) begin
          $fwrite(f, "Register (14,4) Value: %h\n", GRF14_4_buffer[clk]);
        end
        if (GRF14_5_buffer[clk] != GRF14_5_buffer[!clk]) begin
          $fwrite(f, "Register (14,5) Value: %h\n", GRF14_5_buffer[clk]);
        end
        if (GRF14_6_buffer[clk] != GRF14_6_buffer[!clk]) begin
          $fwrite(f, "Register (14,6) Value: %h\n", GRF14_6_buffer[clk]);
        end
        if (GRF14_7_buffer[clk] != GRF14_7_buffer[!clk]) begin
          $fwrite(f, "Register (14,7) Value: %h\n", GRF14_7_buffer[clk]);
        end
        if (GRF14_8_buffer[clk] != GRF14_8_buffer[!clk]) begin
          $fwrite(f, "Register (14,8) Value: %h\n", GRF14_8_buffer[clk]);
        end
        if (GRF14_9_buffer[clk] != GRF14_9_buffer[!clk]) begin
          $fwrite(f, "Register (14,9) Value: %h\n", GRF14_9_buffer[clk]);
        end
        if (GRF14_10_buffer[clk] != GRF14_10_buffer[!clk]) begin
          $fwrite(f, "Register (14,10) Value: %h\n", GRF14_10_buffer[clk]);
        end
        if (GRF14_11_buffer[clk] != GRF14_11_buffer[!clk]) begin
          $fwrite(f, "Register (14,11) Value: %h\n", GRF14_11_buffer[clk]);
        end
        if (GRF14_12_buffer[clk] != GRF14_12_buffer[!clk]) begin
          $fwrite(f, "Register (14,12) Value: %h\n", GRF14_12_buffer[clk]);
        end
        if (GRF14_13_buffer[clk] != GRF14_13_buffer[!clk]) begin
          $fwrite(f, "Register (14,13) Value: %h\n", GRF14_13_buffer[clk]);
        end
        if (GRF14_14_buffer[clk] != GRF14_14_buffer[!clk]) begin
          $fwrite(f, "Register (14,14) Value: %h\n", GRF14_14_buffer[clk]);
        end
        if (GRF14_15_buffer[clk] != GRF14_15_buffer[!clk]) begin
          $fwrite(f, "Register (14,15) Value: %h\n", GRF14_15_buffer[clk]);
        end
        if (GRF14_16_buffer[clk] != GRF14_16_buffer[!clk]) begin
          $fwrite(f, "Register (14,16) Value: %h\n", GRF14_16_buffer[clk]);
        end
        if (GRF14_17_buffer[clk] != GRF14_17_buffer[!clk]) begin
          $fwrite(f, "Register (14,17) Value: %h\n", GRF14_17_buffer[clk]);
        end
        if (GRF14_18_buffer[clk] != GRF14_18_buffer[!clk]) begin
          $fwrite(f, "Register (14,18) Value: %h\n", GRF14_18_buffer[clk]);
        end
        if (GRF14_19_buffer[clk] != GRF14_19_buffer[!clk]) begin
          $fwrite(f, "Register (14,19) Value: %h\n", GRF14_19_buffer[clk]);
        end
        if (GRF14_20_buffer[clk] != GRF14_20_buffer[!clk]) begin
          $fwrite(f, "Register (14,20) Value: %h\n", GRF14_20_buffer[clk]);
        end
        if (GRF14_21_buffer[clk] != GRF14_21_buffer[!clk]) begin
          $fwrite(f, "Register (14,21) Value: %h\n", GRF14_21_buffer[clk]);
        end
        if (GRF14_22_buffer[clk] != GRF14_22_buffer[!clk]) begin
          $fwrite(f, "Register (14,22) Value: %h\n", GRF14_22_buffer[clk]);
        end
        if (GRF14_23_buffer[clk] != GRF14_23_buffer[!clk]) begin
          $fwrite(f, "Register (14,23) Value: %h\n", GRF14_23_buffer[clk]);
        end
        if (GRF14_24_buffer[clk] != GRF14_24_buffer[!clk]) begin
          $fwrite(f, "Register (14,24) Value: %h\n", GRF14_24_buffer[clk]);
        end
        if (GRF14_25_buffer[clk] != GRF14_25_buffer[!clk]) begin
          $fwrite(f, "Register (14,25) Value: %h\n", GRF14_25_buffer[clk]);
        end
        if (GRF14_26_buffer[clk] != GRF14_26_buffer[!clk]) begin
          $fwrite(f, "Register (14,26) Value: %h\n", GRF14_26_buffer[clk]);
        end
        if (GRF14_27_buffer[clk] != GRF14_27_buffer[!clk]) begin
          $fwrite(f, "Register (14,27) Value: %h\n", GRF14_27_buffer[clk]);
        end
        if (GRF14_28_buffer[clk] != GRF14_28_buffer[!clk]) begin
          $fwrite(f, "Register (14,28) Value: %h\n", GRF14_28_buffer[clk]);
        end
        if (GRF14_29_buffer[clk] != GRF14_29_buffer[!clk]) begin
          $fwrite(f, "Register (14,29) Value: %h\n", GRF14_29_buffer[clk]);
        end
        if (GRF14_30_buffer[clk] != GRF14_30_buffer[!clk]) begin
          $fwrite(f, "Register (14,30) Value: %h\n", GRF14_30_buffer[clk]);
        end
        if (GRF14_31_buffer[clk] != GRF14_31_buffer[!clk]) begin
          $fwrite(f, "Register (14,31) Value: %h\n", GRF14_31_buffer[clk]);
        end
        if (GRF15_0_buffer[clk] != GRF15_0_buffer[!clk]) begin
          $fwrite(f, "Register (15,0) Value: %h\n", GRF15_0_buffer[clk]);
        end
        if (GRF15_1_buffer[clk] != GRF15_1_buffer[!clk]) begin
          $fwrite(f, "Register (15,1) Value: %h\n", GRF15_1_buffer[clk]);
        end
        if (GRF15_2_buffer[clk] != GRF15_2_buffer[!clk]) begin
          $fwrite(f, "Register (15,2) Value: %h\n", GRF15_2_buffer[clk]);
        end
        if (GRF15_3_buffer[clk] != GRF15_3_buffer[!clk]) begin
          $fwrite(f, "Register (15,3) Value: %h\n", GRF15_3_buffer[clk]);
        end
        if (GRF15_4_buffer[clk] != GRF15_4_buffer[!clk]) begin
          $fwrite(f, "Register (15,4) Value: %h\n", GRF15_4_buffer[clk]);
        end
        if (GRF15_5_buffer[clk] != GRF15_5_buffer[!clk]) begin
          $fwrite(f, "Register (15,5) Value: %h\n", GRF15_5_buffer[clk]);
        end
        if (GRF15_6_buffer[clk] != GRF15_6_buffer[!clk]) begin
          $fwrite(f, "Register (15,6) Value: %h\n", GRF15_6_buffer[clk]);
        end
        if (GRF15_7_buffer[clk] != GRF15_7_buffer[!clk]) begin
          $fwrite(f, "Register (15,7) Value: %h\n", GRF15_7_buffer[clk]);
        end
        if (GRF15_8_buffer[clk] != GRF15_8_buffer[!clk]) begin
          $fwrite(f, "Register (15,8) Value: %h\n", GRF15_8_buffer[clk]);
        end
        if (GRF15_9_buffer[clk] != GRF15_9_buffer[!clk]) begin
          $fwrite(f, "Register (15,9) Value: %h\n", GRF15_9_buffer[clk]);
        end
        if (GRF15_10_buffer[clk] != GRF15_10_buffer[!clk]) begin
          $fwrite(f, "Register (15,10) Value: %h\n", GRF15_10_buffer[clk]);
        end
        if (GRF15_11_buffer[clk] != GRF15_11_buffer[!clk]) begin
          $fwrite(f, "Register (15,11) Value: %h\n", GRF15_11_buffer[clk]);
        end
        if (GRF15_12_buffer[clk] != GRF15_12_buffer[!clk]) begin
          $fwrite(f, "Register (15,12) Value: %h\n", GRF15_12_buffer[clk]);
        end
        if (GRF15_13_buffer[clk] != GRF15_13_buffer[!clk]) begin
          $fwrite(f, "Register (15,13) Value: %h\n", GRF15_13_buffer[clk]);
        end
        if (GRF15_14_buffer[clk] != GRF15_14_buffer[!clk]) begin
          $fwrite(f, "Register (15,14) Value: %h\n", GRF15_14_buffer[clk]);
        end
        if (GRF15_15_buffer[clk] != GRF15_15_buffer[!clk]) begin
          $fwrite(f, "Register (15,15) Value: %h\n", GRF15_15_buffer[clk]);
        end
        if (GRF15_16_buffer[clk] != GRF15_16_buffer[!clk]) begin
          $fwrite(f, "Register (15,16) Value: %h\n", GRF15_16_buffer[clk]);
        end
        if (GRF15_17_buffer[clk] != GRF15_17_buffer[!clk]) begin
          $fwrite(f, "Register (15,17) Value: %h\n", GRF15_17_buffer[clk]);
        end
        if (GRF15_18_buffer[clk] != GRF15_18_buffer[!clk]) begin
          $fwrite(f, "Register (15,18) Value: %h\n", GRF15_18_buffer[clk]);
        end
        if (GRF15_19_buffer[clk] != GRF15_19_buffer[!clk]) begin
          $fwrite(f, "Register (15,19) Value: %h\n", GRF15_19_buffer[clk]);
        end
        if (GRF15_20_buffer[clk] != GRF15_20_buffer[!clk]) begin
          $fwrite(f, "Register (15,20) Value: %h\n", GRF15_20_buffer[clk]);
        end
        if (GRF15_21_buffer[clk] != GRF15_21_buffer[!clk]) begin
          $fwrite(f, "Register (15,21) Value: %h\n", GRF15_21_buffer[clk]);
        end
        if (GRF15_22_buffer[clk] != GRF15_22_buffer[!clk]) begin
          $fwrite(f, "Register (15,22) Value: %h\n", GRF15_22_buffer[clk]);
        end
        if (GRF15_23_buffer[clk] != GRF15_23_buffer[!clk]) begin
          $fwrite(f, "Register (15,23) Value: %h\n", GRF15_23_buffer[clk]);
        end
        if (GRF15_24_buffer[clk] != GRF15_24_buffer[!clk]) begin
          $fwrite(f, "Register (15,24) Value: %h\n", GRF15_24_buffer[clk]);
        end
        if (GRF15_25_buffer[clk] != GRF15_25_buffer[!clk]) begin
          $fwrite(f, "Register (15,25) Value: %h\n", GRF15_25_buffer[clk]);
        end
        if (GRF15_26_buffer[clk] != GRF15_26_buffer[!clk]) begin
          $fwrite(f, "Register (15,26) Value: %h\n", GRF15_26_buffer[clk]);
        end
        if (GRF15_27_buffer[clk] != GRF15_27_buffer[!clk]) begin
          $fwrite(f, "Register (15,27) Value: %h\n", GRF15_27_buffer[clk]);
        end
        if (GRF15_28_buffer[clk] != GRF15_28_buffer[!clk]) begin
          $fwrite(f, "Register (15,28) Value: %h\n", GRF15_28_buffer[clk]);
        end
        if (GRF15_29_buffer[clk] != GRF15_29_buffer[!clk]) begin
          $fwrite(f, "Register (15,29) Value: %h\n", GRF15_29_buffer[clk]);
        end
        if (GRF15_30_buffer[clk] != GRF15_30_buffer[!clk]) begin
          $fwrite(f, "Register (15,30) Value: %h\n", GRF15_30_buffer[clk]);
        end
        if (GRF15_31_buffer[clk] != GRF15_31_buffer[!clk]) begin
          $fwrite(f, "Register (15,31) Value: %h\n", GRF15_31_buffer[clk]);
        end
        if (GRF16_0_buffer[clk] != GRF16_0_buffer[!clk]) begin
          $fwrite(f, "Register (16,0) Value: %h\n", GRF16_0_buffer[clk]);
        end
        if (GRF16_1_buffer[clk] != GRF16_1_buffer[!clk]) begin
          $fwrite(f, "Register (16,1) Value: %h\n", GRF16_1_buffer[clk]);
        end
        if (GRF16_2_buffer[clk] != GRF16_2_buffer[!clk]) begin
          $fwrite(f, "Register (16,2) Value: %h\n", GRF16_2_buffer[clk]);
        end
        if (GRF16_3_buffer[clk] != GRF16_3_buffer[!clk]) begin
          $fwrite(f, "Register (16,3) Value: %h\n", GRF16_3_buffer[clk]);
        end
        if (GRF16_4_buffer[clk] != GRF16_4_buffer[!clk]) begin
          $fwrite(f, "Register (16,4) Value: %h\n", GRF16_4_buffer[clk]);
        end
        if (GRF16_5_buffer[clk] != GRF16_5_buffer[!clk]) begin
          $fwrite(f, "Register (16,5) Value: %h\n", GRF16_5_buffer[clk]);
        end
        if (GRF16_6_buffer[clk] != GRF16_6_buffer[!clk]) begin
          $fwrite(f, "Register (16,6) Value: %h\n", GRF16_6_buffer[clk]);
        end
        if (GRF16_7_buffer[clk] != GRF16_7_buffer[!clk]) begin
          $fwrite(f, "Register (16,7) Value: %h\n", GRF16_7_buffer[clk]);
        end
        if (GRF16_8_buffer[clk] != GRF16_8_buffer[!clk]) begin
          $fwrite(f, "Register (16,8) Value: %h\n", GRF16_8_buffer[clk]);
        end
        if (GRF16_9_buffer[clk] != GRF16_9_buffer[!clk]) begin
          $fwrite(f, "Register (16,9) Value: %h\n", GRF16_9_buffer[clk]);
        end
        if (GRF16_10_buffer[clk] != GRF16_10_buffer[!clk]) begin
          $fwrite(f, "Register (16,10) Value: %h\n", GRF16_10_buffer[clk]);
        end
        if (GRF16_11_buffer[clk] != GRF16_11_buffer[!clk]) begin
          $fwrite(f, "Register (16,11) Value: %h\n", GRF16_11_buffer[clk]);
        end
        if (GRF16_12_buffer[clk] != GRF16_12_buffer[!clk]) begin
          $fwrite(f, "Register (16,12) Value: %h\n", GRF16_12_buffer[clk]);
        end
        if (GRF16_13_buffer[clk] != GRF16_13_buffer[!clk]) begin
          $fwrite(f, "Register (16,13) Value: %h\n", GRF16_13_buffer[clk]);
        end
        if (GRF16_14_buffer[clk] != GRF16_14_buffer[!clk]) begin
          $fwrite(f, "Register (16,14) Value: %h\n", GRF16_14_buffer[clk]);
        end
        if (GRF16_15_buffer[clk] != GRF16_15_buffer[!clk]) begin
          $fwrite(f, "Register (16,15) Value: %h\n", GRF16_15_buffer[clk]);
        end
        if (GRF16_16_buffer[clk] != GRF16_16_buffer[!clk]) begin
          $fwrite(f, "Register (16,16) Value: %h\n", GRF16_16_buffer[clk]);
        end
        if (GRF16_17_buffer[clk] != GRF16_17_buffer[!clk]) begin
          $fwrite(f, "Register (16,17) Value: %h\n", GRF16_17_buffer[clk]);
        end
        if (GRF16_18_buffer[clk] != GRF16_18_buffer[!clk]) begin
          $fwrite(f, "Register (16,18) Value: %h\n", GRF16_18_buffer[clk]);
        end
        if (GRF16_19_buffer[clk] != GRF16_19_buffer[!clk]) begin
          $fwrite(f, "Register (16,19) Value: %h\n", GRF16_19_buffer[clk]);
        end
        if (GRF16_20_buffer[clk] != GRF16_20_buffer[!clk]) begin
          $fwrite(f, "Register (16,20) Value: %h\n", GRF16_20_buffer[clk]);
        end
        if (GRF16_21_buffer[clk] != GRF16_21_buffer[!clk]) begin
          $fwrite(f, "Register (16,21) Value: %h\n", GRF16_21_buffer[clk]);
        end
        if (GRF16_22_buffer[clk] != GRF16_22_buffer[!clk]) begin
          $fwrite(f, "Register (16,22) Value: %h\n", GRF16_22_buffer[clk]);
        end
        if (GRF16_23_buffer[clk] != GRF16_23_buffer[!clk]) begin
          $fwrite(f, "Register (16,23) Value: %h\n", GRF16_23_buffer[clk]);
        end
        if (GRF16_24_buffer[clk] != GRF16_24_buffer[!clk]) begin
          $fwrite(f, "Register (16,24) Value: %h\n", GRF16_24_buffer[clk]);
        end
        if (GRF16_25_buffer[clk] != GRF16_25_buffer[!clk]) begin
          $fwrite(f, "Register (16,25) Value: %h\n", GRF16_25_buffer[clk]);
        end
        if (GRF16_26_buffer[clk] != GRF16_26_buffer[!clk]) begin
          $fwrite(f, "Register (16,26) Value: %h\n", GRF16_26_buffer[clk]);
        end
        if (GRF16_27_buffer[clk] != GRF16_27_buffer[!clk]) begin
          $fwrite(f, "Register (16,27) Value: %h\n", GRF16_27_buffer[clk]);
        end
        if (GRF16_28_buffer[clk] != GRF16_28_buffer[!clk]) begin
          $fwrite(f, "Register (16,28) Value: %h\n", GRF16_28_buffer[clk]);
        end
        if (GRF16_29_buffer[clk] != GRF16_29_buffer[!clk]) begin
          $fwrite(f, "Register (16,29) Value: %h\n", GRF16_29_buffer[clk]);
        end
        if (GRF16_30_buffer[clk] != GRF16_30_buffer[!clk]) begin
          $fwrite(f, "Register (16,30) Value: %h\n", GRF16_30_buffer[clk]);
        end
        if (GRF16_31_buffer[clk] != GRF16_31_buffer[!clk]) begin
          $fwrite(f, "Register (16,31) Value: %h\n", GRF16_31_buffer[clk]);
        end
        if (GRF17_0_buffer[clk] != GRF17_0_buffer[!clk]) begin
          $fwrite(f, "Register (17,0) Value: %h\n", GRF17_0_buffer[clk]);
        end
        if (GRF17_1_buffer[clk] != GRF17_1_buffer[!clk]) begin
          $fwrite(f, "Register (17,1) Value: %h\n", GRF17_1_buffer[clk]);
        end
        if (GRF17_2_buffer[clk] != GRF17_2_buffer[!clk]) begin
          $fwrite(f, "Register (17,2) Value: %h\n", GRF17_2_buffer[clk]);
        end
        if (GRF17_3_buffer[clk] != GRF17_3_buffer[!clk]) begin
          $fwrite(f, "Register (17,3) Value: %h\n", GRF17_3_buffer[clk]);
        end
        if (GRF17_4_buffer[clk] != GRF17_4_buffer[!clk]) begin
          $fwrite(f, "Register (17,4) Value: %h\n", GRF17_4_buffer[clk]);
        end
        if (GRF17_5_buffer[clk] != GRF17_5_buffer[!clk]) begin
          $fwrite(f, "Register (17,5) Value: %h\n", GRF17_5_buffer[clk]);
        end
        if (GRF17_6_buffer[clk] != GRF17_6_buffer[!clk]) begin
          $fwrite(f, "Register (17,6) Value: %h\n", GRF17_6_buffer[clk]);
        end
        if (GRF17_7_buffer[clk] != GRF17_7_buffer[!clk]) begin
          $fwrite(f, "Register (17,7) Value: %h\n", GRF17_7_buffer[clk]);
        end
        if (GRF17_8_buffer[clk] != GRF17_8_buffer[!clk]) begin
          $fwrite(f, "Register (17,8) Value: %h\n", GRF17_8_buffer[clk]);
        end
        if (GRF17_9_buffer[clk] != GRF17_9_buffer[!clk]) begin
          $fwrite(f, "Register (17,9) Value: %h\n", GRF17_9_buffer[clk]);
        end
        if (GRF17_10_buffer[clk] != GRF17_10_buffer[!clk]) begin
          $fwrite(f, "Register (17,10) Value: %h\n", GRF17_10_buffer[clk]);
        end
        if (GRF17_11_buffer[clk] != GRF17_11_buffer[!clk]) begin
          $fwrite(f, "Register (17,11) Value: %h\n", GRF17_11_buffer[clk]);
        end
        if (GRF17_12_buffer[clk] != GRF17_12_buffer[!clk]) begin
          $fwrite(f, "Register (17,12) Value: %h\n", GRF17_12_buffer[clk]);
        end
        if (GRF17_13_buffer[clk] != GRF17_13_buffer[!clk]) begin
          $fwrite(f, "Register (17,13) Value: %h\n", GRF17_13_buffer[clk]);
        end
        if (GRF17_14_buffer[clk] != GRF17_14_buffer[!clk]) begin
          $fwrite(f, "Register (17,14) Value: %h\n", GRF17_14_buffer[clk]);
        end
        if (GRF17_15_buffer[clk] != GRF17_15_buffer[!clk]) begin
          $fwrite(f, "Register (17,15) Value: %h\n", GRF17_15_buffer[clk]);
        end
        if (GRF17_16_buffer[clk] != GRF17_16_buffer[!clk]) begin
          $fwrite(f, "Register (17,16) Value: %h\n", GRF17_16_buffer[clk]);
        end
        if (GRF17_17_buffer[clk] != GRF17_17_buffer[!clk]) begin
          $fwrite(f, "Register (17,17) Value: %h\n", GRF17_17_buffer[clk]);
        end
        if (GRF17_18_buffer[clk] != GRF17_18_buffer[!clk]) begin
          $fwrite(f, "Register (17,18) Value: %h\n", GRF17_18_buffer[clk]);
        end
        if (GRF17_19_buffer[clk] != GRF17_19_buffer[!clk]) begin
          $fwrite(f, "Register (17,19) Value: %h\n", GRF17_19_buffer[clk]);
        end
        if (GRF17_20_buffer[clk] != GRF17_20_buffer[!clk]) begin
          $fwrite(f, "Register (17,20) Value: %h\n", GRF17_20_buffer[clk]);
        end
        if (GRF17_21_buffer[clk] != GRF17_21_buffer[!clk]) begin
          $fwrite(f, "Register (17,21) Value: %h\n", GRF17_21_buffer[clk]);
        end
        if (GRF17_22_buffer[clk] != GRF17_22_buffer[!clk]) begin
          $fwrite(f, "Register (17,22) Value: %h\n", GRF17_22_buffer[clk]);
        end
        if (GRF17_23_buffer[clk] != GRF17_23_buffer[!clk]) begin
          $fwrite(f, "Register (17,23) Value: %h\n", GRF17_23_buffer[clk]);
        end
        if (GRF17_24_buffer[clk] != GRF17_24_buffer[!clk]) begin
          $fwrite(f, "Register (17,24) Value: %h\n", GRF17_24_buffer[clk]);
        end
        if (GRF17_25_buffer[clk] != GRF17_25_buffer[!clk]) begin
          $fwrite(f, "Register (17,25) Value: %h\n", GRF17_25_buffer[clk]);
        end
        if (GRF17_26_buffer[clk] != GRF17_26_buffer[!clk]) begin
          $fwrite(f, "Register (17,26) Value: %h\n", GRF17_26_buffer[clk]);
        end
        if (GRF17_27_buffer[clk] != GRF17_27_buffer[!clk]) begin
          $fwrite(f, "Register (17,27) Value: %h\n", GRF17_27_buffer[clk]);
        end
        if (GRF17_28_buffer[clk] != GRF17_28_buffer[!clk]) begin
          $fwrite(f, "Register (17,28) Value: %h\n", GRF17_28_buffer[clk]);
        end
        if (GRF17_29_buffer[clk] != GRF17_29_buffer[!clk]) begin
          $fwrite(f, "Register (17,29) Value: %h\n", GRF17_29_buffer[clk]);
        end
        if (GRF17_30_buffer[clk] != GRF17_30_buffer[!clk]) begin
          $fwrite(f, "Register (17,30) Value: %h\n", GRF17_30_buffer[clk]);
        end
        if (GRF17_31_buffer[clk] != GRF17_31_buffer[!clk]) begin
          $fwrite(f, "Register (17,31) Value: %h\n", GRF17_31_buffer[clk]);
        end
        if (GRF18_0_buffer[clk] != GRF18_0_buffer[!clk]) begin
          $fwrite(f, "Register (18,0) Value: %h\n", GRF18_0_buffer[clk]);
        end
        if (GRF18_1_buffer[clk] != GRF18_1_buffer[!clk]) begin
          $fwrite(f, "Register (18,1) Value: %h\n", GRF18_1_buffer[clk]);
        end
        if (GRF18_2_buffer[clk] != GRF18_2_buffer[!clk]) begin
          $fwrite(f, "Register (18,2) Value: %h\n", GRF18_2_buffer[clk]);
        end
        if (GRF18_3_buffer[clk] != GRF18_3_buffer[!clk]) begin
          $fwrite(f, "Register (18,3) Value: %h\n", GRF18_3_buffer[clk]);
        end
        if (GRF18_4_buffer[clk] != GRF18_4_buffer[!clk]) begin
          $fwrite(f, "Register (18,4) Value: %h\n", GRF18_4_buffer[clk]);
        end
        if (GRF18_5_buffer[clk] != GRF18_5_buffer[!clk]) begin
          $fwrite(f, "Register (18,5) Value: %h\n", GRF18_5_buffer[clk]);
        end
        if (GRF18_6_buffer[clk] != GRF18_6_buffer[!clk]) begin
          $fwrite(f, "Register (18,6) Value: %h\n", GRF18_6_buffer[clk]);
        end
        if (GRF18_7_buffer[clk] != GRF18_7_buffer[!clk]) begin
          $fwrite(f, "Register (18,7) Value: %h\n", GRF18_7_buffer[clk]);
        end
        if (GRF18_8_buffer[clk] != GRF18_8_buffer[!clk]) begin
          $fwrite(f, "Register (18,8) Value: %h\n", GRF18_8_buffer[clk]);
        end
        if (GRF18_9_buffer[clk] != GRF18_9_buffer[!clk]) begin
          $fwrite(f, "Register (18,9) Value: %h\n", GRF18_9_buffer[clk]);
        end
        if (GRF18_10_buffer[clk] != GRF18_10_buffer[!clk]) begin
          $fwrite(f, "Register (18,10) Value: %h\n", GRF18_10_buffer[clk]);
        end
        if (GRF18_11_buffer[clk] != GRF18_11_buffer[!clk]) begin
          $fwrite(f, "Register (18,11) Value: %h\n", GRF18_11_buffer[clk]);
        end
        if (GRF18_12_buffer[clk] != GRF18_12_buffer[!clk]) begin
          $fwrite(f, "Register (18,12) Value: %h\n", GRF18_12_buffer[clk]);
        end
        if (GRF18_13_buffer[clk] != GRF18_13_buffer[!clk]) begin
          $fwrite(f, "Register (18,13) Value: %h\n", GRF18_13_buffer[clk]);
        end
        if (GRF18_14_buffer[clk] != GRF18_14_buffer[!clk]) begin
          $fwrite(f, "Register (18,14) Value: %h\n", GRF18_14_buffer[clk]);
        end
        if (GRF18_15_buffer[clk] != GRF18_15_buffer[!clk]) begin
          $fwrite(f, "Register (18,15) Value: %h\n", GRF18_15_buffer[clk]);
        end
        if (GRF18_16_buffer[clk] != GRF18_16_buffer[!clk]) begin
          $fwrite(f, "Register (18,16) Value: %h\n", GRF18_16_buffer[clk]);
        end
        if (GRF18_17_buffer[clk] != GRF18_17_buffer[!clk]) begin
          $fwrite(f, "Register (18,17) Value: %h\n", GRF18_17_buffer[clk]);
        end
        if (GRF18_18_buffer[clk] != GRF18_18_buffer[!clk]) begin
          $fwrite(f, "Register (18,18) Value: %h\n", GRF18_18_buffer[clk]);
        end
        if (GRF18_19_buffer[clk] != GRF18_19_buffer[!clk]) begin
          $fwrite(f, "Register (18,19) Value: %h\n", GRF18_19_buffer[clk]);
        end
        if (GRF18_20_buffer[clk] != GRF18_20_buffer[!clk]) begin
          $fwrite(f, "Register (18,20) Value: %h\n", GRF18_20_buffer[clk]);
        end
        if (GRF18_21_buffer[clk] != GRF18_21_buffer[!clk]) begin
          $fwrite(f, "Register (18,21) Value: %h\n", GRF18_21_buffer[clk]);
        end
        if (GRF18_22_buffer[clk] != GRF18_22_buffer[!clk]) begin
          $fwrite(f, "Register (18,22) Value: %h\n", GRF18_22_buffer[clk]);
        end
        if (GRF18_23_buffer[clk] != GRF18_23_buffer[!clk]) begin
          $fwrite(f, "Register (18,23) Value: %h\n", GRF18_23_buffer[clk]);
        end
        if (GRF18_24_buffer[clk] != GRF18_24_buffer[!clk]) begin
          $fwrite(f, "Register (18,24) Value: %h\n", GRF18_24_buffer[clk]);
        end
        if (GRF18_25_buffer[clk] != GRF18_25_buffer[!clk]) begin
          $fwrite(f, "Register (18,25) Value: %h\n", GRF18_25_buffer[clk]);
        end
        if (GRF18_26_buffer[clk] != GRF18_26_buffer[!clk]) begin
          $fwrite(f, "Register (18,26) Value: %h\n", GRF18_26_buffer[clk]);
        end
        if (GRF18_27_buffer[clk] != GRF18_27_buffer[!clk]) begin
          $fwrite(f, "Register (18,27) Value: %h\n", GRF18_27_buffer[clk]);
        end
        if (GRF18_28_buffer[clk] != GRF18_28_buffer[!clk]) begin
          $fwrite(f, "Register (18,28) Value: %h\n", GRF18_28_buffer[clk]);
        end
        if (GRF18_29_buffer[clk] != GRF18_29_buffer[!clk]) begin
          $fwrite(f, "Register (18,29) Value: %h\n", GRF18_29_buffer[clk]);
        end
        if (GRF18_30_buffer[clk] != GRF18_30_buffer[!clk]) begin
          $fwrite(f, "Register (18,30) Value: %h\n", GRF18_30_buffer[clk]);
        end
        if (GRF18_31_buffer[clk] != GRF18_31_buffer[!clk]) begin
          $fwrite(f, "Register (18,31) Value: %h\n", GRF18_31_buffer[clk]);
        end
        if (GRF19_0_buffer[clk] != GRF19_0_buffer[!clk]) begin
          $fwrite(f, "Register (19,0) Value: %h\n", GRF19_0_buffer[clk]);
        end
        if (GRF19_1_buffer[clk] != GRF19_1_buffer[!clk]) begin
          $fwrite(f, "Register (19,1) Value: %h\n", GRF19_1_buffer[clk]);
        end
        if (GRF19_2_buffer[clk] != GRF19_2_buffer[!clk]) begin
          $fwrite(f, "Register (19,2) Value: %h\n", GRF19_2_buffer[clk]);
        end
        if (GRF19_3_buffer[clk] != GRF19_3_buffer[!clk]) begin
          $fwrite(f, "Register (19,3) Value: %h\n", GRF19_3_buffer[clk]);
        end
        if (GRF19_4_buffer[clk] != GRF19_4_buffer[!clk]) begin
          $fwrite(f, "Register (19,4) Value: %h\n", GRF19_4_buffer[clk]);
        end
        if (GRF19_5_buffer[clk] != GRF19_5_buffer[!clk]) begin
          $fwrite(f, "Register (19,5) Value: %h\n", GRF19_5_buffer[clk]);
        end
        if (GRF19_6_buffer[clk] != GRF19_6_buffer[!clk]) begin
          $fwrite(f, "Register (19,6) Value: %h\n", GRF19_6_buffer[clk]);
        end
        if (GRF19_7_buffer[clk] != GRF19_7_buffer[!clk]) begin
          $fwrite(f, "Register (19,7) Value: %h\n", GRF19_7_buffer[clk]);
        end
        if (GRF19_8_buffer[clk] != GRF19_8_buffer[!clk]) begin
          $fwrite(f, "Register (19,8) Value: %h\n", GRF19_8_buffer[clk]);
        end
        if (GRF19_9_buffer[clk] != GRF19_9_buffer[!clk]) begin
          $fwrite(f, "Register (19,9) Value: %h\n", GRF19_9_buffer[clk]);
        end
        if (GRF19_10_buffer[clk] != GRF19_10_buffer[!clk]) begin
          $fwrite(f, "Register (19,10) Value: %h\n", GRF19_10_buffer[clk]);
        end
        if (GRF19_11_buffer[clk] != GRF19_11_buffer[!clk]) begin
          $fwrite(f, "Register (19,11) Value: %h\n", GRF19_11_buffer[clk]);
        end
        if (GRF19_12_buffer[clk] != GRF19_12_buffer[!clk]) begin
          $fwrite(f, "Register (19,12) Value: %h\n", GRF19_12_buffer[clk]);
        end
        if (GRF19_13_buffer[clk] != GRF19_13_buffer[!clk]) begin
          $fwrite(f, "Register (19,13) Value: %h\n", GRF19_13_buffer[clk]);
        end
        if (GRF19_14_buffer[clk] != GRF19_14_buffer[!clk]) begin
          $fwrite(f, "Register (19,14) Value: %h\n", GRF19_14_buffer[clk]);
        end
        if (GRF19_15_buffer[clk] != GRF19_15_buffer[!clk]) begin
          $fwrite(f, "Register (19,15) Value: %h\n", GRF19_15_buffer[clk]);
        end
        if (GRF19_16_buffer[clk] != GRF19_16_buffer[!clk]) begin
          $fwrite(f, "Register (19,16) Value: %h\n", GRF19_16_buffer[clk]);
        end
        if (GRF19_17_buffer[clk] != GRF19_17_buffer[!clk]) begin
          $fwrite(f, "Register (19,17) Value: %h\n", GRF19_17_buffer[clk]);
        end
        if (GRF19_18_buffer[clk] != GRF19_18_buffer[!clk]) begin
          $fwrite(f, "Register (19,18) Value: %h\n", GRF19_18_buffer[clk]);
        end
        if (GRF19_19_buffer[clk] != GRF19_19_buffer[!clk]) begin
          $fwrite(f, "Register (19,19) Value: %h\n", GRF19_19_buffer[clk]);
        end
        if (GRF19_20_buffer[clk] != GRF19_20_buffer[!clk]) begin
          $fwrite(f, "Register (19,20) Value: %h\n", GRF19_20_buffer[clk]);
        end
        if (GRF19_21_buffer[clk] != GRF19_21_buffer[!clk]) begin
          $fwrite(f, "Register (19,21) Value: %h\n", GRF19_21_buffer[clk]);
        end
        if (GRF19_22_buffer[clk] != GRF19_22_buffer[!clk]) begin
          $fwrite(f, "Register (19,22) Value: %h\n", GRF19_22_buffer[clk]);
        end
        if (GRF19_23_buffer[clk] != GRF19_23_buffer[!clk]) begin
          $fwrite(f, "Register (19,23) Value: %h\n", GRF19_23_buffer[clk]);
        end
        if (GRF19_24_buffer[clk] != GRF19_24_buffer[!clk]) begin
          $fwrite(f, "Register (19,24) Value: %h\n", GRF19_24_buffer[clk]);
        end
        if (GRF19_25_buffer[clk] != GRF19_25_buffer[!clk]) begin
          $fwrite(f, "Register (19,25) Value: %h\n", GRF19_25_buffer[clk]);
        end
        if (GRF19_26_buffer[clk] != GRF19_26_buffer[!clk]) begin
          $fwrite(f, "Register (19,26) Value: %h\n", GRF19_26_buffer[clk]);
        end
        if (GRF19_27_buffer[clk] != GRF19_27_buffer[!clk]) begin
          $fwrite(f, "Register (19,27) Value: %h\n", GRF19_27_buffer[clk]);
        end
        if (GRF19_28_buffer[clk] != GRF19_28_buffer[!clk]) begin
          $fwrite(f, "Register (19,28) Value: %h\n", GRF19_28_buffer[clk]);
        end
        if (GRF19_29_buffer[clk] != GRF19_29_buffer[!clk]) begin
          $fwrite(f, "Register (19,29) Value: %h\n", GRF19_29_buffer[clk]);
        end
        if (GRF19_30_buffer[clk] != GRF19_30_buffer[!clk]) begin
          $fwrite(f, "Register (19,30) Value: %h\n", GRF19_30_buffer[clk]);
        end
        if (GRF19_31_buffer[clk] != GRF19_31_buffer[!clk]) begin
          $fwrite(f, "Register (19,31) Value: %h\n", GRF19_31_buffer[clk]);
        end
        if (GRF20_0_buffer[clk] != GRF20_0_buffer[!clk]) begin
          $fwrite(f, "Register (20,0) Value: %h\n", GRF20_0_buffer[clk]);
        end
        if (GRF20_1_buffer[clk] != GRF20_1_buffer[!clk]) begin
          $fwrite(f, "Register (20,1) Value: %h\n", GRF20_1_buffer[clk]);
        end
        if (GRF20_2_buffer[clk] != GRF20_2_buffer[!clk]) begin
          $fwrite(f, "Register (20,2) Value: %h\n", GRF20_2_buffer[clk]);
        end
        if (GRF20_3_buffer[clk] != GRF20_3_buffer[!clk]) begin
          $fwrite(f, "Register (20,3) Value: %h\n", GRF20_3_buffer[clk]);
        end
        if (GRF20_4_buffer[clk] != GRF20_4_buffer[!clk]) begin
          $fwrite(f, "Register (20,4) Value: %h\n", GRF20_4_buffer[clk]);
        end
        if (GRF20_5_buffer[clk] != GRF20_5_buffer[!clk]) begin
          $fwrite(f, "Register (20,5) Value: %h\n", GRF20_5_buffer[clk]);
        end
        if (GRF20_6_buffer[clk] != GRF20_6_buffer[!clk]) begin
          $fwrite(f, "Register (20,6) Value: %h\n", GRF20_6_buffer[clk]);
        end
        if (GRF20_7_buffer[clk] != GRF20_7_buffer[!clk]) begin
          $fwrite(f, "Register (20,7) Value: %h\n", GRF20_7_buffer[clk]);
        end
        if (GRF20_8_buffer[clk] != GRF20_8_buffer[!clk]) begin
          $fwrite(f, "Register (20,8) Value: %h\n", GRF20_8_buffer[clk]);
        end
        if (GRF20_9_buffer[clk] != GRF20_9_buffer[!clk]) begin
          $fwrite(f, "Register (20,9) Value: %h\n", GRF20_9_buffer[clk]);
        end
        if (GRF20_10_buffer[clk] != GRF20_10_buffer[!clk]) begin
          $fwrite(f, "Register (20,10) Value: %h\n", GRF20_10_buffer[clk]);
        end
        if (GRF20_11_buffer[clk] != GRF20_11_buffer[!clk]) begin
          $fwrite(f, "Register (20,11) Value: %h\n", GRF20_11_buffer[clk]);
        end
        if (GRF20_12_buffer[clk] != GRF20_12_buffer[!clk]) begin
          $fwrite(f, "Register (20,12) Value: %h\n", GRF20_12_buffer[clk]);
        end
        if (GRF20_13_buffer[clk] != GRF20_13_buffer[!clk]) begin
          $fwrite(f, "Register (20,13) Value: %h\n", GRF20_13_buffer[clk]);
        end
        if (GRF20_14_buffer[clk] != GRF20_14_buffer[!clk]) begin
          $fwrite(f, "Register (20,14) Value: %h\n", GRF20_14_buffer[clk]);
        end
        if (GRF20_15_buffer[clk] != GRF20_15_buffer[!clk]) begin
          $fwrite(f, "Register (20,15) Value: %h\n", GRF20_15_buffer[clk]);
        end
        if (GRF20_16_buffer[clk] != GRF20_16_buffer[!clk]) begin
          $fwrite(f, "Register (20,16) Value: %h\n", GRF20_16_buffer[clk]);
        end
        if (GRF20_17_buffer[clk] != GRF20_17_buffer[!clk]) begin
          $fwrite(f, "Register (20,17) Value: %h\n", GRF20_17_buffer[clk]);
        end
        if (GRF20_18_buffer[clk] != GRF20_18_buffer[!clk]) begin
          $fwrite(f, "Register (20,18) Value: %h\n", GRF20_18_buffer[clk]);
        end
        if (GRF20_19_buffer[clk] != GRF20_19_buffer[!clk]) begin
          $fwrite(f, "Register (20,19) Value: %h\n", GRF20_19_buffer[clk]);
        end
        if (GRF20_20_buffer[clk] != GRF20_20_buffer[!clk]) begin
          $fwrite(f, "Register (20,20) Value: %h\n", GRF20_20_buffer[clk]);
        end
        if (GRF20_21_buffer[clk] != GRF20_21_buffer[!clk]) begin
          $fwrite(f, "Register (20,21) Value: %h\n", GRF20_21_buffer[clk]);
        end
        if (GRF20_22_buffer[clk] != GRF20_22_buffer[!clk]) begin
          $fwrite(f, "Register (20,22) Value: %h\n", GRF20_22_buffer[clk]);
        end
        if (GRF20_23_buffer[clk] != GRF20_23_buffer[!clk]) begin
          $fwrite(f, "Register (20,23) Value: %h\n", GRF20_23_buffer[clk]);
        end
        if (GRF20_24_buffer[clk] != GRF20_24_buffer[!clk]) begin
          $fwrite(f, "Register (20,24) Value: %h\n", GRF20_24_buffer[clk]);
        end
        if (GRF20_25_buffer[clk] != GRF20_25_buffer[!clk]) begin
          $fwrite(f, "Register (20,25) Value: %h\n", GRF20_25_buffer[clk]);
        end
        if (GRF20_26_buffer[clk] != GRF20_26_buffer[!clk]) begin
          $fwrite(f, "Register (20,26) Value: %h\n", GRF20_26_buffer[clk]);
        end
        if (GRF20_27_buffer[clk] != GRF20_27_buffer[!clk]) begin
          $fwrite(f, "Register (20,27) Value: %h\n", GRF20_27_buffer[clk]);
        end
        if (GRF20_28_buffer[clk] != GRF20_28_buffer[!clk]) begin
          $fwrite(f, "Register (20,28) Value: %h\n", GRF20_28_buffer[clk]);
        end
        if (GRF20_29_buffer[clk] != GRF20_29_buffer[!clk]) begin
          $fwrite(f, "Register (20,29) Value: %h\n", GRF20_29_buffer[clk]);
        end
        if (GRF20_30_buffer[clk] != GRF20_30_buffer[!clk]) begin
          $fwrite(f, "Register (20,30) Value: %h\n", GRF20_30_buffer[clk]);
        end
        if (GRF20_31_buffer[clk] != GRF20_31_buffer[!clk]) begin
          $fwrite(f, "Register (20,31) Value: %h\n", GRF20_31_buffer[clk]);
        end
        if (GRF21_0_buffer[clk] != GRF21_0_buffer[!clk]) begin
          $fwrite(f, "Register (21,0) Value: %h\n", GRF21_0_buffer[clk]);
        end
        if (GRF21_1_buffer[clk] != GRF21_1_buffer[!clk]) begin
          $fwrite(f, "Register (21,1) Value: %h\n", GRF21_1_buffer[clk]);
        end
        if (GRF21_2_buffer[clk] != GRF21_2_buffer[!clk]) begin
          $fwrite(f, "Register (21,2) Value: %h\n", GRF21_2_buffer[clk]);
        end
        if (GRF21_3_buffer[clk] != GRF21_3_buffer[!clk]) begin
          $fwrite(f, "Register (21,3) Value: %h\n", GRF21_3_buffer[clk]);
        end
        if (GRF21_4_buffer[clk] != GRF21_4_buffer[!clk]) begin
          $fwrite(f, "Register (21,4) Value: %h\n", GRF21_4_buffer[clk]);
        end
        if (GRF21_5_buffer[clk] != GRF21_5_buffer[!clk]) begin
          $fwrite(f, "Register (21,5) Value: %h\n", GRF21_5_buffer[clk]);
        end
        if (GRF21_6_buffer[clk] != GRF21_6_buffer[!clk]) begin
          $fwrite(f, "Register (21,6) Value: %h\n", GRF21_6_buffer[clk]);
        end
        if (GRF21_7_buffer[clk] != GRF21_7_buffer[!clk]) begin
          $fwrite(f, "Register (21,7) Value: %h\n", GRF21_7_buffer[clk]);
        end
        if (GRF21_8_buffer[clk] != GRF21_8_buffer[!clk]) begin
          $fwrite(f, "Register (21,8) Value: %h\n", GRF21_8_buffer[clk]);
        end
        if (GRF21_9_buffer[clk] != GRF21_9_buffer[!clk]) begin
          $fwrite(f, "Register (21,9) Value: %h\n", GRF21_9_buffer[clk]);
        end
        if (GRF21_10_buffer[clk] != GRF21_10_buffer[!clk]) begin
          $fwrite(f, "Register (21,10) Value: %h\n", GRF21_10_buffer[clk]);
        end
        if (GRF21_11_buffer[clk] != GRF21_11_buffer[!clk]) begin
          $fwrite(f, "Register (21,11) Value: %h\n", GRF21_11_buffer[clk]);
        end
        if (GRF21_12_buffer[clk] != GRF21_12_buffer[!clk]) begin
          $fwrite(f, "Register (21,12) Value: %h\n", GRF21_12_buffer[clk]);
        end
        if (GRF21_13_buffer[clk] != GRF21_13_buffer[!clk]) begin
          $fwrite(f, "Register (21,13) Value: %h\n", GRF21_13_buffer[clk]);
        end
        if (GRF21_14_buffer[clk] != GRF21_14_buffer[!clk]) begin
          $fwrite(f, "Register (21,14) Value: %h\n", GRF21_14_buffer[clk]);
        end
        if (GRF21_15_buffer[clk] != GRF21_15_buffer[!clk]) begin
          $fwrite(f, "Register (21,15) Value: %h\n", GRF21_15_buffer[clk]);
        end
        if (GRF21_16_buffer[clk] != GRF21_16_buffer[!clk]) begin
          $fwrite(f, "Register (21,16) Value: %h\n", GRF21_16_buffer[clk]);
        end
        if (GRF21_17_buffer[clk] != GRF21_17_buffer[!clk]) begin
          $fwrite(f, "Register (21,17) Value: %h\n", GRF21_17_buffer[clk]);
        end
        if (GRF21_18_buffer[clk] != GRF21_18_buffer[!clk]) begin
          $fwrite(f, "Register (21,18) Value: %h\n", GRF21_18_buffer[clk]);
        end
        if (GRF21_19_buffer[clk] != GRF21_19_buffer[!clk]) begin
          $fwrite(f, "Register (21,19) Value: %h\n", GRF21_19_buffer[clk]);
        end
        if (GRF21_20_buffer[clk] != GRF21_20_buffer[!clk]) begin
          $fwrite(f, "Register (21,20) Value: %h\n", GRF21_20_buffer[clk]);
        end
        if (GRF21_21_buffer[clk] != GRF21_21_buffer[!clk]) begin
          $fwrite(f, "Register (21,21) Value: %h\n", GRF21_21_buffer[clk]);
        end
        if (GRF21_22_buffer[clk] != GRF21_22_buffer[!clk]) begin
          $fwrite(f, "Register (21,22) Value: %h\n", GRF21_22_buffer[clk]);
        end
        if (GRF21_23_buffer[clk] != GRF21_23_buffer[!clk]) begin
          $fwrite(f, "Register (21,23) Value: %h\n", GRF21_23_buffer[clk]);
        end
        if (GRF21_24_buffer[clk] != GRF21_24_buffer[!clk]) begin
          $fwrite(f, "Register (21,24) Value: %h\n", GRF21_24_buffer[clk]);
        end
        if (GRF21_25_buffer[clk] != GRF21_25_buffer[!clk]) begin
          $fwrite(f, "Register (21,25) Value: %h\n", GRF21_25_buffer[clk]);
        end
        if (GRF21_26_buffer[clk] != GRF21_26_buffer[!clk]) begin
          $fwrite(f, "Register (21,26) Value: %h\n", GRF21_26_buffer[clk]);
        end
        if (GRF21_27_buffer[clk] != GRF21_27_buffer[!clk]) begin
          $fwrite(f, "Register (21,27) Value: %h\n", GRF21_27_buffer[clk]);
        end
        if (GRF21_28_buffer[clk] != GRF21_28_buffer[!clk]) begin
          $fwrite(f, "Register (21,28) Value: %h\n", GRF21_28_buffer[clk]);
        end
        if (GRF21_29_buffer[clk] != GRF21_29_buffer[!clk]) begin
          $fwrite(f, "Register (21,29) Value: %h\n", GRF21_29_buffer[clk]);
        end
        if (GRF21_30_buffer[clk] != GRF21_30_buffer[!clk]) begin
          $fwrite(f, "Register (21,30) Value: %h\n", GRF21_30_buffer[clk]);
        end
        if (GRF21_31_buffer[clk] != GRF21_31_buffer[!clk]) begin
          $fwrite(f, "Register (21,31) Value: %h\n", GRF21_31_buffer[clk]);
        end
        if (GRF22_0_buffer[clk] != GRF22_0_buffer[!clk]) begin
          $fwrite(f, "Register (22,0) Value: %h\n", GRF22_0_buffer[clk]);
        end
        if (GRF22_1_buffer[clk] != GRF22_1_buffer[!clk]) begin
          $fwrite(f, "Register (22,1) Value: %h\n", GRF22_1_buffer[clk]);
        end
        if (GRF22_2_buffer[clk] != GRF22_2_buffer[!clk]) begin
          $fwrite(f, "Register (22,2) Value: %h\n", GRF22_2_buffer[clk]);
        end
        if (GRF22_3_buffer[clk] != GRF22_3_buffer[!clk]) begin
          $fwrite(f, "Register (22,3) Value: %h\n", GRF22_3_buffer[clk]);
        end
        if (GRF22_4_buffer[clk] != GRF22_4_buffer[!clk]) begin
          $fwrite(f, "Register (22,4) Value: %h\n", GRF22_4_buffer[clk]);
        end
        if (GRF22_5_buffer[clk] != GRF22_5_buffer[!clk]) begin
          $fwrite(f, "Register (22,5) Value: %h\n", GRF22_5_buffer[clk]);
        end
        if (GRF22_6_buffer[clk] != GRF22_6_buffer[!clk]) begin
          $fwrite(f, "Register (22,6) Value: %h\n", GRF22_6_buffer[clk]);
        end
        if (GRF22_7_buffer[clk] != GRF22_7_buffer[!clk]) begin
          $fwrite(f, "Register (22,7) Value: %h\n", GRF22_7_buffer[clk]);
        end
        if (GRF22_8_buffer[clk] != GRF22_8_buffer[!clk]) begin
          $fwrite(f, "Register (22,8) Value: %h\n", GRF22_8_buffer[clk]);
        end
        if (GRF22_9_buffer[clk] != GRF22_9_buffer[!clk]) begin
          $fwrite(f, "Register (22,9) Value: %h\n", GRF22_9_buffer[clk]);
        end
        if (GRF22_10_buffer[clk] != GRF22_10_buffer[!clk]) begin
          $fwrite(f, "Register (22,10) Value: %h\n", GRF22_10_buffer[clk]);
        end
        if (GRF22_11_buffer[clk] != GRF22_11_buffer[!clk]) begin
          $fwrite(f, "Register (22,11) Value: %h\n", GRF22_11_buffer[clk]);
        end
        if (GRF22_12_buffer[clk] != GRF22_12_buffer[!clk]) begin
          $fwrite(f, "Register (22,12) Value: %h\n", GRF22_12_buffer[clk]);
        end
        if (GRF22_13_buffer[clk] != GRF22_13_buffer[!clk]) begin
          $fwrite(f, "Register (22,13) Value: %h\n", GRF22_13_buffer[clk]);
        end
        if (GRF22_14_buffer[clk] != GRF22_14_buffer[!clk]) begin
          $fwrite(f, "Register (22,14) Value: %h\n", GRF22_14_buffer[clk]);
        end
        if (GRF22_15_buffer[clk] != GRF22_15_buffer[!clk]) begin
          $fwrite(f, "Register (22,15) Value: %h\n", GRF22_15_buffer[clk]);
        end
        if (GRF22_16_buffer[clk] != GRF22_16_buffer[!clk]) begin
          $fwrite(f, "Register (22,16) Value: %h\n", GRF22_16_buffer[clk]);
        end
        if (GRF22_17_buffer[clk] != GRF22_17_buffer[!clk]) begin
          $fwrite(f, "Register (22,17) Value: %h\n", GRF22_17_buffer[clk]);
        end
        if (GRF22_18_buffer[clk] != GRF22_18_buffer[!clk]) begin
          $fwrite(f, "Register (22,18) Value: %h\n", GRF22_18_buffer[clk]);
        end
        if (GRF22_19_buffer[clk] != GRF22_19_buffer[!clk]) begin
          $fwrite(f, "Register (22,19) Value: %h\n", GRF22_19_buffer[clk]);
        end
        if (GRF22_20_buffer[clk] != GRF22_20_buffer[!clk]) begin
          $fwrite(f, "Register (22,20) Value: %h\n", GRF22_20_buffer[clk]);
        end
        if (GRF22_21_buffer[clk] != GRF22_21_buffer[!clk]) begin
          $fwrite(f, "Register (22,21) Value: %h\n", GRF22_21_buffer[clk]);
        end
        if (GRF22_22_buffer[clk] != GRF22_22_buffer[!clk]) begin
          $fwrite(f, "Register (22,22) Value: %h\n", GRF22_22_buffer[clk]);
        end
        if (GRF22_23_buffer[clk] != GRF22_23_buffer[!clk]) begin
          $fwrite(f, "Register (22,23) Value: %h\n", GRF22_23_buffer[clk]);
        end
        if (GRF22_24_buffer[clk] != GRF22_24_buffer[!clk]) begin
          $fwrite(f, "Register (22,24) Value: %h\n", GRF22_24_buffer[clk]);
        end
        if (GRF22_25_buffer[clk] != GRF22_25_buffer[!clk]) begin
          $fwrite(f, "Register (22,25) Value: %h\n", GRF22_25_buffer[clk]);
        end
        if (GRF22_26_buffer[clk] != GRF22_26_buffer[!clk]) begin
          $fwrite(f, "Register (22,26) Value: %h\n", GRF22_26_buffer[clk]);
        end
        if (GRF22_27_buffer[clk] != GRF22_27_buffer[!clk]) begin
          $fwrite(f, "Register (22,27) Value: %h\n", GRF22_27_buffer[clk]);
        end
        if (GRF22_28_buffer[clk] != GRF22_28_buffer[!clk]) begin
          $fwrite(f, "Register (22,28) Value: %h\n", GRF22_28_buffer[clk]);
        end
        if (GRF22_29_buffer[clk] != GRF22_29_buffer[!clk]) begin
          $fwrite(f, "Register (22,29) Value: %h\n", GRF22_29_buffer[clk]);
        end
        if (GRF22_30_buffer[clk] != GRF22_30_buffer[!clk]) begin
          $fwrite(f, "Register (22,30) Value: %h\n", GRF22_30_buffer[clk]);
        end
        if (GRF22_31_buffer[clk] != GRF22_31_buffer[!clk]) begin
          $fwrite(f, "Register (22,31) Value: %h\n", GRF22_31_buffer[clk]);
        end
        if (GRF23_0_buffer[clk] != GRF23_0_buffer[!clk]) begin
          $fwrite(f, "Register (23,0) Value: %h\n", GRF23_0_buffer[clk]);
        end
        if (GRF23_1_buffer[clk] != GRF23_1_buffer[!clk]) begin
          $fwrite(f, "Register (23,1) Value: %h\n", GRF23_1_buffer[clk]);
        end
        if (GRF23_2_buffer[clk] != GRF23_2_buffer[!clk]) begin
          $fwrite(f, "Register (23,2) Value: %h\n", GRF23_2_buffer[clk]);
        end
        if (GRF23_3_buffer[clk] != GRF23_3_buffer[!clk]) begin
          $fwrite(f, "Register (23,3) Value: %h\n", GRF23_3_buffer[clk]);
        end
        if (GRF23_4_buffer[clk] != GRF23_4_buffer[!clk]) begin
          $fwrite(f, "Register (23,4) Value: %h\n", GRF23_4_buffer[clk]);
        end
        if (GRF23_5_buffer[clk] != GRF23_5_buffer[!clk]) begin
          $fwrite(f, "Register (23,5) Value: %h\n", GRF23_5_buffer[clk]);
        end
        if (GRF23_6_buffer[clk] != GRF23_6_buffer[!clk]) begin
          $fwrite(f, "Register (23,6) Value: %h\n", GRF23_6_buffer[clk]);
        end
        if (GRF23_7_buffer[clk] != GRF23_7_buffer[!clk]) begin
          $fwrite(f, "Register (23,7) Value: %h\n", GRF23_7_buffer[clk]);
        end
        if (GRF23_8_buffer[clk] != GRF23_8_buffer[!clk]) begin
          $fwrite(f, "Register (23,8) Value: %h\n", GRF23_8_buffer[clk]);
        end
        if (GRF23_9_buffer[clk] != GRF23_9_buffer[!clk]) begin
          $fwrite(f, "Register (23,9) Value: %h\n", GRF23_9_buffer[clk]);
        end
        if (GRF23_10_buffer[clk] != GRF23_10_buffer[!clk]) begin
          $fwrite(f, "Register (23,10) Value: %h\n", GRF23_10_buffer[clk]);
        end
        if (GRF23_11_buffer[clk] != GRF23_11_buffer[!clk]) begin
          $fwrite(f, "Register (23,11) Value: %h\n", GRF23_11_buffer[clk]);
        end
        if (GRF23_12_buffer[clk] != GRF23_12_buffer[!clk]) begin
          $fwrite(f, "Register (23,12) Value: %h\n", GRF23_12_buffer[clk]);
        end
        if (GRF23_13_buffer[clk] != GRF23_13_buffer[!clk]) begin
          $fwrite(f, "Register (23,13) Value: %h\n", GRF23_13_buffer[clk]);
        end
        if (GRF23_14_buffer[clk] != GRF23_14_buffer[!clk]) begin
          $fwrite(f, "Register (23,14) Value: %h\n", GRF23_14_buffer[clk]);
        end
        if (GRF23_15_buffer[clk] != GRF23_15_buffer[!clk]) begin
          $fwrite(f, "Register (23,15) Value: %h\n", GRF23_15_buffer[clk]);
        end
        if (GRF23_16_buffer[clk] != GRF23_16_buffer[!clk]) begin
          $fwrite(f, "Register (23,16) Value: %h\n", GRF23_16_buffer[clk]);
        end
        if (GRF23_17_buffer[clk] != GRF23_17_buffer[!clk]) begin
          $fwrite(f, "Register (23,17) Value: %h\n", GRF23_17_buffer[clk]);
        end
        if (GRF23_18_buffer[clk] != GRF23_18_buffer[!clk]) begin
          $fwrite(f, "Register (23,18) Value: %h\n", GRF23_18_buffer[clk]);
        end
        if (GRF23_19_buffer[clk] != GRF23_19_buffer[!clk]) begin
          $fwrite(f, "Register (23,19) Value: %h\n", GRF23_19_buffer[clk]);
        end
        if (GRF23_20_buffer[clk] != GRF23_20_buffer[!clk]) begin
          $fwrite(f, "Register (23,20) Value: %h\n", GRF23_20_buffer[clk]);
        end
        if (GRF23_21_buffer[clk] != GRF23_21_buffer[!clk]) begin
          $fwrite(f, "Register (23,21) Value: %h\n", GRF23_21_buffer[clk]);
        end
        if (GRF23_22_buffer[clk] != GRF23_22_buffer[!clk]) begin
          $fwrite(f, "Register (23,22) Value: %h\n", GRF23_22_buffer[clk]);
        end
        if (GRF23_23_buffer[clk] != GRF23_23_buffer[!clk]) begin
          $fwrite(f, "Register (23,23) Value: %h\n", GRF23_23_buffer[clk]);
        end
        if (GRF23_24_buffer[clk] != GRF23_24_buffer[!clk]) begin
          $fwrite(f, "Register (23,24) Value: %h\n", GRF23_24_buffer[clk]);
        end
        if (GRF23_25_buffer[clk] != GRF23_25_buffer[!clk]) begin
          $fwrite(f, "Register (23,25) Value: %h\n", GRF23_25_buffer[clk]);
        end
        if (GRF23_26_buffer[clk] != GRF23_26_buffer[!clk]) begin
          $fwrite(f, "Register (23,26) Value: %h\n", GRF23_26_buffer[clk]);
        end
        if (GRF23_27_buffer[clk] != GRF23_27_buffer[!clk]) begin
          $fwrite(f, "Register (23,27) Value: %h\n", GRF23_27_buffer[clk]);
        end
        if (GRF23_28_buffer[clk] != GRF23_28_buffer[!clk]) begin
          $fwrite(f, "Register (23,28) Value: %h\n", GRF23_28_buffer[clk]);
        end
        if (GRF23_29_buffer[clk] != GRF23_29_buffer[!clk]) begin
          $fwrite(f, "Register (23,29) Value: %h\n", GRF23_29_buffer[clk]);
        end
        if (GRF23_30_buffer[clk] != GRF23_30_buffer[!clk]) begin
          $fwrite(f, "Register (23,30) Value: %h\n", GRF23_30_buffer[clk]);
        end
        if (GRF23_31_buffer[clk] != GRF23_31_buffer[!clk]) begin
          $fwrite(f, "Register (23,31) Value: %h\n", GRF23_31_buffer[clk]);
        end
        if (GRF24_0_buffer[clk] != GRF24_0_buffer[!clk]) begin
          $fwrite(f, "Register (24,0) Value: %h\n", GRF24_0_buffer[clk]);
        end
        if (GRF24_1_buffer[clk] != GRF24_1_buffer[!clk]) begin
          $fwrite(f, "Register (24,1) Value: %h\n", GRF24_1_buffer[clk]);
        end
        if (GRF24_2_buffer[clk] != GRF24_2_buffer[!clk]) begin
          $fwrite(f, "Register (24,2) Value: %h\n", GRF24_2_buffer[clk]);
        end
        if (GRF24_3_buffer[clk] != GRF24_3_buffer[!clk]) begin
          $fwrite(f, "Register (24,3) Value: %h\n", GRF24_3_buffer[clk]);
        end
        if (GRF24_4_buffer[clk] != GRF24_4_buffer[!clk]) begin
          $fwrite(f, "Register (24,4) Value: %h\n", GRF24_4_buffer[clk]);
        end
        if (GRF24_5_buffer[clk] != GRF24_5_buffer[!clk]) begin
          $fwrite(f, "Register (24,5) Value: %h\n", GRF24_5_buffer[clk]);
        end
        if (GRF24_6_buffer[clk] != GRF24_6_buffer[!clk]) begin
          $fwrite(f, "Register (24,6) Value: %h\n", GRF24_6_buffer[clk]);
        end
        if (GRF24_7_buffer[clk] != GRF24_7_buffer[!clk]) begin
          $fwrite(f, "Register (24,7) Value: %h\n", GRF24_7_buffer[clk]);
        end
        if (GRF24_8_buffer[clk] != GRF24_8_buffer[!clk]) begin
          $fwrite(f, "Register (24,8) Value: %h\n", GRF24_8_buffer[clk]);
        end
        if (GRF24_9_buffer[clk] != GRF24_9_buffer[!clk]) begin
          $fwrite(f, "Register (24,9) Value: %h\n", GRF24_9_buffer[clk]);
        end
        if (GRF24_10_buffer[clk] != GRF24_10_buffer[!clk]) begin
          $fwrite(f, "Register (24,10) Value: %h\n", GRF24_10_buffer[clk]);
        end
        if (GRF24_11_buffer[clk] != GRF24_11_buffer[!clk]) begin
          $fwrite(f, "Register (24,11) Value: %h\n", GRF24_11_buffer[clk]);
        end
        if (GRF24_12_buffer[clk] != GRF24_12_buffer[!clk]) begin
          $fwrite(f, "Register (24,12) Value: %h\n", GRF24_12_buffer[clk]);
        end
        if (GRF24_13_buffer[clk] != GRF24_13_buffer[!clk]) begin
          $fwrite(f, "Register (24,13) Value: %h\n", GRF24_13_buffer[clk]);
        end
        if (GRF24_14_buffer[clk] != GRF24_14_buffer[!clk]) begin
          $fwrite(f, "Register (24,14) Value: %h\n", GRF24_14_buffer[clk]);
        end
        if (GRF24_15_buffer[clk] != GRF24_15_buffer[!clk]) begin
          $fwrite(f, "Register (24,15) Value: %h\n", GRF24_15_buffer[clk]);
        end
        if (GRF24_16_buffer[clk] != GRF24_16_buffer[!clk]) begin
          $fwrite(f, "Register (24,16) Value: %h\n", GRF24_16_buffer[clk]);
        end
        if (GRF24_17_buffer[clk] != GRF24_17_buffer[!clk]) begin
          $fwrite(f, "Register (24,17) Value: %h\n", GRF24_17_buffer[clk]);
        end
        if (GRF24_18_buffer[clk] != GRF24_18_buffer[!clk]) begin
          $fwrite(f, "Register (24,18) Value: %h\n", GRF24_18_buffer[clk]);
        end
        if (GRF24_19_buffer[clk] != GRF24_19_buffer[!clk]) begin
          $fwrite(f, "Register (24,19) Value: %h\n", GRF24_19_buffer[clk]);
        end
        if (GRF24_20_buffer[clk] != GRF24_20_buffer[!clk]) begin
          $fwrite(f, "Register (24,20) Value: %h\n", GRF24_20_buffer[clk]);
        end
        if (GRF24_21_buffer[clk] != GRF24_21_buffer[!clk]) begin
          $fwrite(f, "Register (24,21) Value: %h\n", GRF24_21_buffer[clk]);
        end
        if (GRF24_22_buffer[clk] != GRF24_22_buffer[!clk]) begin
          $fwrite(f, "Register (24,22) Value: %h\n", GRF24_22_buffer[clk]);
        end
        if (GRF24_23_buffer[clk] != GRF24_23_buffer[!clk]) begin
          $fwrite(f, "Register (24,23) Value: %h\n", GRF24_23_buffer[clk]);
        end
        if (GRF24_24_buffer[clk] != GRF24_24_buffer[!clk]) begin
          $fwrite(f, "Register (24,24) Value: %h\n", GRF24_24_buffer[clk]);
        end
        if (GRF24_25_buffer[clk] != GRF24_25_buffer[!clk]) begin
          $fwrite(f, "Register (24,25) Value: %h\n", GRF24_25_buffer[clk]);
        end
        if (GRF24_26_buffer[clk] != GRF24_26_buffer[!clk]) begin
          $fwrite(f, "Register (24,26) Value: %h\n", GRF24_26_buffer[clk]);
        end
        if (GRF24_27_buffer[clk] != GRF24_27_buffer[!clk]) begin
          $fwrite(f, "Register (24,27) Value: %h\n", GRF24_27_buffer[clk]);
        end
        if (GRF24_28_buffer[clk] != GRF24_28_buffer[!clk]) begin
          $fwrite(f, "Register (24,28) Value: %h\n", GRF24_28_buffer[clk]);
        end
        if (GRF24_29_buffer[clk] != GRF24_29_buffer[!clk]) begin
          $fwrite(f, "Register (24,29) Value: %h\n", GRF24_29_buffer[clk]);
        end
        if (GRF24_30_buffer[clk] != GRF24_30_buffer[!clk]) begin
          $fwrite(f, "Register (24,30) Value: %h\n", GRF24_30_buffer[clk]);
        end
        if (GRF24_31_buffer[clk] != GRF24_31_buffer[!clk]) begin
          $fwrite(f, "Register (24,31) Value: %h\n", GRF24_31_buffer[clk]);
        end
        if (GRF25_0_buffer[clk] != GRF25_0_buffer[!clk]) begin
          $fwrite(f, "Register (25,0) Value: %h\n", GRF25_0_buffer[clk]);
        end
        if (GRF25_1_buffer[clk] != GRF25_1_buffer[!clk]) begin
          $fwrite(f, "Register (25,1) Value: %h\n", GRF25_1_buffer[clk]);
        end
        if (GRF25_2_buffer[clk] != GRF25_2_buffer[!clk]) begin
          $fwrite(f, "Register (25,2) Value: %h\n", GRF25_2_buffer[clk]);
        end
        if (GRF25_3_buffer[clk] != GRF25_3_buffer[!clk]) begin
          $fwrite(f, "Register (25,3) Value: %h\n", GRF25_3_buffer[clk]);
        end
        if (GRF25_4_buffer[clk] != GRF25_4_buffer[!clk]) begin
          $fwrite(f, "Register (25,4) Value: %h\n", GRF25_4_buffer[clk]);
        end
        if (GRF25_5_buffer[clk] != GRF25_5_buffer[!clk]) begin
          $fwrite(f, "Register (25,5) Value: %h\n", GRF25_5_buffer[clk]);
        end
        if (GRF25_6_buffer[clk] != GRF25_6_buffer[!clk]) begin
          $fwrite(f, "Register (25,6) Value: %h\n", GRF25_6_buffer[clk]);
        end
        if (GRF25_7_buffer[clk] != GRF25_7_buffer[!clk]) begin
          $fwrite(f, "Register (25,7) Value: %h\n", GRF25_7_buffer[clk]);
        end
        if (GRF25_8_buffer[clk] != GRF25_8_buffer[!clk]) begin
          $fwrite(f, "Register (25,8) Value: %h\n", GRF25_8_buffer[clk]);
        end
        if (GRF25_9_buffer[clk] != GRF25_9_buffer[!clk]) begin
          $fwrite(f, "Register (25,9) Value: %h\n", GRF25_9_buffer[clk]);
        end
        if (GRF25_10_buffer[clk] != GRF25_10_buffer[!clk]) begin
          $fwrite(f, "Register (25,10) Value: %h\n", GRF25_10_buffer[clk]);
        end
        if (GRF25_11_buffer[clk] != GRF25_11_buffer[!clk]) begin
          $fwrite(f, "Register (25,11) Value: %h\n", GRF25_11_buffer[clk]);
        end
        if (GRF25_12_buffer[clk] != GRF25_12_buffer[!clk]) begin
          $fwrite(f, "Register (25,12) Value: %h\n", GRF25_12_buffer[clk]);
        end
        if (GRF25_13_buffer[clk] != GRF25_13_buffer[!clk]) begin
          $fwrite(f, "Register (25,13) Value: %h\n", GRF25_13_buffer[clk]);
        end
        if (GRF25_14_buffer[clk] != GRF25_14_buffer[!clk]) begin
          $fwrite(f, "Register (25,14) Value: %h\n", GRF25_14_buffer[clk]);
        end
        if (GRF25_15_buffer[clk] != GRF25_15_buffer[!clk]) begin
          $fwrite(f, "Register (25,15) Value: %h\n", GRF25_15_buffer[clk]);
        end
        if (GRF25_16_buffer[clk] != GRF25_16_buffer[!clk]) begin
          $fwrite(f, "Register (25,16) Value: %h\n", GRF25_16_buffer[clk]);
        end
        if (GRF25_17_buffer[clk] != GRF25_17_buffer[!clk]) begin
          $fwrite(f, "Register (25,17) Value: %h\n", GRF25_17_buffer[clk]);
        end
        if (GRF25_18_buffer[clk] != GRF25_18_buffer[!clk]) begin
          $fwrite(f, "Register (25,18) Value: %h\n", GRF25_18_buffer[clk]);
        end
        if (GRF25_19_buffer[clk] != GRF25_19_buffer[!clk]) begin
          $fwrite(f, "Register (25,19) Value: %h\n", GRF25_19_buffer[clk]);
        end
        if (GRF25_20_buffer[clk] != GRF25_20_buffer[!clk]) begin
          $fwrite(f, "Register (25,20) Value: %h\n", GRF25_20_buffer[clk]);
        end
        if (GRF25_21_buffer[clk] != GRF25_21_buffer[!clk]) begin
          $fwrite(f, "Register (25,21) Value: %h\n", GRF25_21_buffer[clk]);
        end
        if (GRF25_22_buffer[clk] != GRF25_22_buffer[!clk]) begin
          $fwrite(f, "Register (25,22) Value: %h\n", GRF25_22_buffer[clk]);
        end
        if (GRF25_23_buffer[clk] != GRF25_23_buffer[!clk]) begin
          $fwrite(f, "Register (25,23) Value: %h\n", GRF25_23_buffer[clk]);
        end
        if (GRF25_24_buffer[clk] != GRF25_24_buffer[!clk]) begin
          $fwrite(f, "Register (25,24) Value: %h\n", GRF25_24_buffer[clk]);
        end
        if (GRF25_25_buffer[clk] != GRF25_25_buffer[!clk]) begin
          $fwrite(f, "Register (25,25) Value: %h\n", GRF25_25_buffer[clk]);
        end
        if (GRF25_26_buffer[clk] != GRF25_26_buffer[!clk]) begin
          $fwrite(f, "Register (25,26) Value: %h\n", GRF25_26_buffer[clk]);
        end
        if (GRF25_27_buffer[clk] != GRF25_27_buffer[!clk]) begin
          $fwrite(f, "Register (25,27) Value: %h\n", GRF25_27_buffer[clk]);
        end
        if (GRF25_28_buffer[clk] != GRF25_28_buffer[!clk]) begin
          $fwrite(f, "Register (25,28) Value: %h\n", GRF25_28_buffer[clk]);
        end
        if (GRF25_29_buffer[clk] != GRF25_29_buffer[!clk]) begin
          $fwrite(f, "Register (25,29) Value: %h\n", GRF25_29_buffer[clk]);
        end
        if (GRF25_30_buffer[clk] != GRF25_30_buffer[!clk]) begin
          $fwrite(f, "Register (25,30) Value: %h\n", GRF25_30_buffer[clk]);
        end
        if (GRF25_31_buffer[clk] != GRF25_31_buffer[!clk]) begin
          $fwrite(f, "Register (25,31) Value: %h\n", GRF25_31_buffer[clk]);
        end
        if (GRF26_0_buffer[clk] != GRF26_0_buffer[!clk]) begin
          $fwrite(f, "Register (26,0) Value: %h\n", GRF26_0_buffer[clk]);
        end
        if (GRF26_1_buffer[clk] != GRF26_1_buffer[!clk]) begin
          $fwrite(f, "Register (26,1) Value: %h\n", GRF26_1_buffer[clk]);
        end
        if (GRF26_2_buffer[clk] != GRF26_2_buffer[!clk]) begin
          $fwrite(f, "Register (26,2) Value: %h\n", GRF26_2_buffer[clk]);
        end
        if (GRF26_3_buffer[clk] != GRF26_3_buffer[!clk]) begin
          $fwrite(f, "Register (26,3) Value: %h\n", GRF26_3_buffer[clk]);
        end
        if (GRF26_4_buffer[clk] != GRF26_4_buffer[!clk]) begin
          $fwrite(f, "Register (26,4) Value: %h\n", GRF26_4_buffer[clk]);
        end
        if (GRF26_5_buffer[clk] != GRF26_5_buffer[!clk]) begin
          $fwrite(f, "Register (26,5) Value: %h\n", GRF26_5_buffer[clk]);
        end
        if (GRF26_6_buffer[clk] != GRF26_6_buffer[!clk]) begin
          $fwrite(f, "Register (26,6) Value: %h\n", GRF26_6_buffer[clk]);
        end
        if (GRF26_7_buffer[clk] != GRF26_7_buffer[!clk]) begin
          $fwrite(f, "Register (26,7) Value: %h\n", GRF26_7_buffer[clk]);
        end
        if (GRF26_8_buffer[clk] != GRF26_8_buffer[!clk]) begin
          $fwrite(f, "Register (26,8) Value: %h\n", GRF26_8_buffer[clk]);
        end
        if (GRF26_9_buffer[clk] != GRF26_9_buffer[!clk]) begin
          $fwrite(f, "Register (26,9) Value: %h\n", GRF26_9_buffer[clk]);
        end
        if (GRF26_10_buffer[clk] != GRF26_10_buffer[!clk]) begin
          $fwrite(f, "Register (26,10) Value: %h\n", GRF26_10_buffer[clk]);
        end
        if (GRF26_11_buffer[clk] != GRF26_11_buffer[!clk]) begin
          $fwrite(f, "Register (26,11) Value: %h\n", GRF26_11_buffer[clk]);
        end
        if (GRF26_12_buffer[clk] != GRF26_12_buffer[!clk]) begin
          $fwrite(f, "Register (26,12) Value: %h\n", GRF26_12_buffer[clk]);
        end
        if (GRF26_13_buffer[clk] != GRF26_13_buffer[!clk]) begin
          $fwrite(f, "Register (26,13) Value: %h\n", GRF26_13_buffer[clk]);
        end
        if (GRF26_14_buffer[clk] != GRF26_14_buffer[!clk]) begin
          $fwrite(f, "Register (26,14) Value: %h\n", GRF26_14_buffer[clk]);
        end
        if (GRF26_15_buffer[clk] != GRF26_15_buffer[!clk]) begin
          $fwrite(f, "Register (26,15) Value: %h\n", GRF26_15_buffer[clk]);
        end
        if (GRF26_16_buffer[clk] != GRF26_16_buffer[!clk]) begin
          $fwrite(f, "Register (26,16) Value: %h\n", GRF26_16_buffer[clk]);
        end
        if (GRF26_17_buffer[clk] != GRF26_17_buffer[!clk]) begin
          $fwrite(f, "Register (26,17) Value: %h\n", GRF26_17_buffer[clk]);
        end
        if (GRF26_18_buffer[clk] != GRF26_18_buffer[!clk]) begin
          $fwrite(f, "Register (26,18) Value: %h\n", GRF26_18_buffer[clk]);
        end
        if (GRF26_19_buffer[clk] != GRF26_19_buffer[!clk]) begin
          $fwrite(f, "Register (26,19) Value: %h\n", GRF26_19_buffer[clk]);
        end
        if (GRF26_20_buffer[clk] != GRF26_20_buffer[!clk]) begin
          $fwrite(f, "Register (26,20) Value: %h\n", GRF26_20_buffer[clk]);
        end
        if (GRF26_21_buffer[clk] != GRF26_21_buffer[!clk]) begin
          $fwrite(f, "Register (26,21) Value: %h\n", GRF26_21_buffer[clk]);
        end
        if (GRF26_22_buffer[clk] != GRF26_22_buffer[!clk]) begin
          $fwrite(f, "Register (26,22) Value: %h\n", GRF26_22_buffer[clk]);
        end
        if (GRF26_23_buffer[clk] != GRF26_23_buffer[!clk]) begin
          $fwrite(f, "Register (26,23) Value: %h\n", GRF26_23_buffer[clk]);
        end
        if (GRF26_24_buffer[clk] != GRF26_24_buffer[!clk]) begin
          $fwrite(f, "Register (26,24) Value: %h\n", GRF26_24_buffer[clk]);
        end
        if (GRF26_25_buffer[clk] != GRF26_25_buffer[!clk]) begin
          $fwrite(f, "Register (26,25) Value: %h\n", GRF26_25_buffer[clk]);
        end
        if (GRF26_26_buffer[clk] != GRF26_26_buffer[!clk]) begin
          $fwrite(f, "Register (26,26) Value: %h\n", GRF26_26_buffer[clk]);
        end
        if (GRF26_27_buffer[clk] != GRF26_27_buffer[!clk]) begin
          $fwrite(f, "Register (26,27) Value: %h\n", GRF26_27_buffer[clk]);
        end
        if (GRF26_28_buffer[clk] != GRF26_28_buffer[!clk]) begin
          $fwrite(f, "Register (26,28) Value: %h\n", GRF26_28_buffer[clk]);
        end
        if (GRF26_29_buffer[clk] != GRF26_29_buffer[!clk]) begin
          $fwrite(f, "Register (26,29) Value: %h\n", GRF26_29_buffer[clk]);
        end
        if (GRF26_30_buffer[clk] != GRF26_30_buffer[!clk]) begin
          $fwrite(f, "Register (26,30) Value: %h\n", GRF26_30_buffer[clk]);
        end
        if (GRF26_31_buffer[clk] != GRF26_31_buffer[!clk]) begin
          $fwrite(f, "Register (26,31) Value: %h\n", GRF26_31_buffer[clk]);
        end
        if (GRF27_0_buffer[clk] != GRF27_0_buffer[!clk]) begin
          $fwrite(f, "Register (27,0) Value: %h\n", GRF27_0_buffer[clk]);
        end
        if (GRF27_1_buffer[clk] != GRF27_1_buffer[!clk]) begin
          $fwrite(f, "Register (27,1) Value: %h\n", GRF27_1_buffer[clk]);
        end
        if (GRF27_2_buffer[clk] != GRF27_2_buffer[!clk]) begin
          $fwrite(f, "Register (27,2) Value: %h\n", GRF27_2_buffer[clk]);
        end
        if (GRF27_3_buffer[clk] != GRF27_3_buffer[!clk]) begin
          $fwrite(f, "Register (27,3) Value: %h\n", GRF27_3_buffer[clk]);
        end
        if (GRF27_4_buffer[clk] != GRF27_4_buffer[!clk]) begin
          $fwrite(f, "Register (27,4) Value: %h\n", GRF27_4_buffer[clk]);
        end
        if (GRF27_5_buffer[clk] != GRF27_5_buffer[!clk]) begin
          $fwrite(f, "Register (27,5) Value: %h\n", GRF27_5_buffer[clk]);
        end
        if (GRF27_6_buffer[clk] != GRF27_6_buffer[!clk]) begin
          $fwrite(f, "Register (27,6) Value: %h\n", GRF27_6_buffer[clk]);
        end
        if (GRF27_7_buffer[clk] != GRF27_7_buffer[!clk]) begin
          $fwrite(f, "Register (27,7) Value: %h\n", GRF27_7_buffer[clk]);
        end
        if (GRF27_8_buffer[clk] != GRF27_8_buffer[!clk]) begin
          $fwrite(f, "Register (27,8) Value: %h\n", GRF27_8_buffer[clk]);
        end
        if (GRF27_9_buffer[clk] != GRF27_9_buffer[!clk]) begin
          $fwrite(f, "Register (27,9) Value: %h\n", GRF27_9_buffer[clk]);
        end
        if (GRF27_10_buffer[clk] != GRF27_10_buffer[!clk]) begin
          $fwrite(f, "Register (27,10) Value: %h\n", GRF27_10_buffer[clk]);
        end
        if (GRF27_11_buffer[clk] != GRF27_11_buffer[!clk]) begin
          $fwrite(f, "Register (27,11) Value: %h\n", GRF27_11_buffer[clk]);
        end
        if (GRF27_12_buffer[clk] != GRF27_12_buffer[!clk]) begin
          $fwrite(f, "Register (27,12) Value: %h\n", GRF27_12_buffer[clk]);
        end
        if (GRF27_13_buffer[clk] != GRF27_13_buffer[!clk]) begin
          $fwrite(f, "Register (27,13) Value: %h\n", GRF27_13_buffer[clk]);
        end
        if (GRF27_14_buffer[clk] != GRF27_14_buffer[!clk]) begin
          $fwrite(f, "Register (27,14) Value: %h\n", GRF27_14_buffer[clk]);
        end
        if (GRF27_15_buffer[clk] != GRF27_15_buffer[!clk]) begin
          $fwrite(f, "Register (27,15) Value: %h\n", GRF27_15_buffer[clk]);
        end
        if (GRF27_16_buffer[clk] != GRF27_16_buffer[!clk]) begin
          $fwrite(f, "Register (27,16) Value: %h\n", GRF27_16_buffer[clk]);
        end
        if (GRF27_17_buffer[clk] != GRF27_17_buffer[!clk]) begin
          $fwrite(f, "Register (27,17) Value: %h\n", GRF27_17_buffer[clk]);
        end
        if (GRF27_18_buffer[clk] != GRF27_18_buffer[!clk]) begin
          $fwrite(f, "Register (27,18) Value: %h\n", GRF27_18_buffer[clk]);
        end
        if (GRF27_19_buffer[clk] != GRF27_19_buffer[!clk]) begin
          $fwrite(f, "Register (27,19) Value: %h\n", GRF27_19_buffer[clk]);
        end
        if (GRF27_20_buffer[clk] != GRF27_20_buffer[!clk]) begin
          $fwrite(f, "Register (27,20) Value: %h\n", GRF27_20_buffer[clk]);
        end
        if (GRF27_21_buffer[clk] != GRF27_21_buffer[!clk]) begin
          $fwrite(f, "Register (27,21) Value: %h\n", GRF27_21_buffer[clk]);
        end
        if (GRF27_22_buffer[clk] != GRF27_22_buffer[!clk]) begin
          $fwrite(f, "Register (27,22) Value: %h\n", GRF27_22_buffer[clk]);
        end
        if (GRF27_23_buffer[clk] != GRF27_23_buffer[!clk]) begin
          $fwrite(f, "Register (27,23) Value: %h\n", GRF27_23_buffer[clk]);
        end
        if (GRF27_24_buffer[clk] != GRF27_24_buffer[!clk]) begin
          $fwrite(f, "Register (27,24) Value: %h\n", GRF27_24_buffer[clk]);
        end
        if (GRF27_25_buffer[clk] != GRF27_25_buffer[!clk]) begin
          $fwrite(f, "Register (27,25) Value: %h\n", GRF27_25_buffer[clk]);
        end
        if (GRF27_26_buffer[clk] != GRF27_26_buffer[!clk]) begin
          $fwrite(f, "Register (27,26) Value: %h\n", GRF27_26_buffer[clk]);
        end
        if (GRF27_27_buffer[clk] != GRF27_27_buffer[!clk]) begin
          $fwrite(f, "Register (27,27) Value: %h\n", GRF27_27_buffer[clk]);
        end
        if (GRF27_28_buffer[clk] != GRF27_28_buffer[!clk]) begin
          $fwrite(f, "Register (27,28) Value: %h\n", GRF27_28_buffer[clk]);
        end
        if (GRF27_29_buffer[clk] != GRF27_29_buffer[!clk]) begin
          $fwrite(f, "Register (27,29) Value: %h\n", GRF27_29_buffer[clk]);
        end
        if (GRF27_30_buffer[clk] != GRF27_30_buffer[!clk]) begin
          $fwrite(f, "Register (27,30) Value: %h\n", GRF27_30_buffer[clk]);
        end
        if (GRF27_31_buffer[clk] != GRF27_31_buffer[!clk]) begin
          $fwrite(f, "Register (27,31) Value: %h\n", GRF27_31_buffer[clk]);
        end
        if (GRF28_0_buffer[clk] != GRF28_0_buffer[!clk]) begin
          $fwrite(f, "Register (28,0) Value: %h\n", GRF28_0_buffer[clk]);
        end
        if (GRF28_1_buffer[clk] != GRF28_1_buffer[!clk]) begin
          $fwrite(f, "Register (28,1) Value: %h\n", GRF28_1_buffer[clk]);
        end
        if (GRF28_2_buffer[clk] != GRF28_2_buffer[!clk]) begin
          $fwrite(f, "Register (28,2) Value: %h\n", GRF28_2_buffer[clk]);
        end
        if (GRF28_3_buffer[clk] != GRF28_3_buffer[!clk]) begin
          $fwrite(f, "Register (28,3) Value: %h\n", GRF28_3_buffer[clk]);
        end
        if (GRF28_4_buffer[clk] != GRF28_4_buffer[!clk]) begin
          $fwrite(f, "Register (28,4) Value: %h\n", GRF28_4_buffer[clk]);
        end
        if (GRF28_5_buffer[clk] != GRF28_5_buffer[!clk]) begin
          $fwrite(f, "Register (28,5) Value: %h\n", GRF28_5_buffer[clk]);
        end
        if (GRF28_6_buffer[clk] != GRF28_6_buffer[!clk]) begin
          $fwrite(f, "Register (28,6) Value: %h\n", GRF28_6_buffer[clk]);
        end
        if (GRF28_7_buffer[clk] != GRF28_7_buffer[!clk]) begin
          $fwrite(f, "Register (28,7) Value: %h\n", GRF28_7_buffer[clk]);
        end
        if (GRF28_8_buffer[clk] != GRF28_8_buffer[!clk]) begin
          $fwrite(f, "Register (28,8) Value: %h\n", GRF28_8_buffer[clk]);
        end
        if (GRF28_9_buffer[clk] != GRF28_9_buffer[!clk]) begin
          $fwrite(f, "Register (28,9) Value: %h\n", GRF28_9_buffer[clk]);
        end
        if (GRF28_10_buffer[clk] != GRF28_10_buffer[!clk]) begin
          $fwrite(f, "Register (28,10) Value: %h\n", GRF28_10_buffer[clk]);
        end
        if (GRF28_11_buffer[clk] != GRF28_11_buffer[!clk]) begin
          $fwrite(f, "Register (28,11) Value: %h\n", GRF28_11_buffer[clk]);
        end
        if (GRF28_12_buffer[clk] != GRF28_12_buffer[!clk]) begin
          $fwrite(f, "Register (28,12) Value: %h\n", GRF28_12_buffer[clk]);
        end
        if (GRF28_13_buffer[clk] != GRF28_13_buffer[!clk]) begin
          $fwrite(f, "Register (28,13) Value: %h\n", GRF28_13_buffer[clk]);
        end
        if (GRF28_14_buffer[clk] != GRF28_14_buffer[!clk]) begin
          $fwrite(f, "Register (28,14) Value: %h\n", GRF28_14_buffer[clk]);
        end
        if (GRF28_15_buffer[clk] != GRF28_15_buffer[!clk]) begin
          $fwrite(f, "Register (28,15) Value: %h\n", GRF28_15_buffer[clk]);
        end
        if (GRF28_16_buffer[clk] != GRF28_16_buffer[!clk]) begin
          $fwrite(f, "Register (28,16) Value: %h\n", GRF28_16_buffer[clk]);
        end
        if (GRF28_17_buffer[clk] != GRF28_17_buffer[!clk]) begin
          $fwrite(f, "Register (28,17) Value: %h\n", GRF28_17_buffer[clk]);
        end
        if (GRF28_18_buffer[clk] != GRF28_18_buffer[!clk]) begin
          $fwrite(f, "Register (28,18) Value: %h\n", GRF28_18_buffer[clk]);
        end
        if (GRF28_19_buffer[clk] != GRF28_19_buffer[!clk]) begin
          $fwrite(f, "Register (28,19) Value: %h\n", GRF28_19_buffer[clk]);
        end
        if (GRF28_20_buffer[clk] != GRF28_20_buffer[!clk]) begin
          $fwrite(f, "Register (28,20) Value: %h\n", GRF28_20_buffer[clk]);
        end
        if (GRF28_21_buffer[clk] != GRF28_21_buffer[!clk]) begin
          $fwrite(f, "Register (28,21) Value: %h\n", GRF28_21_buffer[clk]);
        end
        if (GRF28_22_buffer[clk] != GRF28_22_buffer[!clk]) begin
          $fwrite(f, "Register (28,22) Value: %h\n", GRF28_22_buffer[clk]);
        end
        if (GRF28_23_buffer[clk] != GRF28_23_buffer[!clk]) begin
          $fwrite(f, "Register (28,23) Value: %h\n", GRF28_23_buffer[clk]);
        end
        if (GRF28_24_buffer[clk] != GRF28_24_buffer[!clk]) begin
          $fwrite(f, "Register (28,24) Value: %h\n", GRF28_24_buffer[clk]);
        end
        if (GRF28_25_buffer[clk] != GRF28_25_buffer[!clk]) begin
          $fwrite(f, "Register (28,25) Value: %h\n", GRF28_25_buffer[clk]);
        end
        if (GRF28_26_buffer[clk] != GRF28_26_buffer[!clk]) begin
          $fwrite(f, "Register (28,26) Value: %h\n", GRF28_26_buffer[clk]);
        end
        if (GRF28_27_buffer[clk] != GRF28_27_buffer[!clk]) begin
          $fwrite(f, "Register (28,27) Value: %h\n", GRF28_27_buffer[clk]);
        end
        if (GRF28_28_buffer[clk] != GRF28_28_buffer[!clk]) begin
          $fwrite(f, "Register (28,28) Value: %h\n", GRF28_28_buffer[clk]);
        end
        if (GRF28_29_buffer[clk] != GRF28_29_buffer[!clk]) begin
          $fwrite(f, "Register (28,29) Value: %h\n", GRF28_29_buffer[clk]);
        end
        if (GRF28_30_buffer[clk] != GRF28_30_buffer[!clk]) begin
          $fwrite(f, "Register (28,30) Value: %h\n", GRF28_30_buffer[clk]);
        end
        if (GRF28_31_buffer[clk] != GRF28_31_buffer[!clk]) begin
          $fwrite(f, "Register (28,31) Value: %h\n", GRF28_31_buffer[clk]);
        end
        if (GRF29_0_buffer[clk] != GRF29_0_buffer[!clk]) begin
          $fwrite(f, "Register (29,0) Value: %h\n", GRF29_0_buffer[clk]);
        end
        if (GRF29_1_buffer[clk] != GRF29_1_buffer[!clk]) begin
          $fwrite(f, "Register (29,1) Value: %h\n", GRF29_1_buffer[clk]);
        end
        if (GRF29_2_buffer[clk] != GRF29_2_buffer[!clk]) begin
          $fwrite(f, "Register (29,2) Value: %h\n", GRF29_2_buffer[clk]);
        end
        if (GRF29_3_buffer[clk] != GRF29_3_buffer[!clk]) begin
          $fwrite(f, "Register (29,3) Value: %h\n", GRF29_3_buffer[clk]);
        end
        if (GRF29_4_buffer[clk] != GRF29_4_buffer[!clk]) begin
          $fwrite(f, "Register (29,4) Value: %h\n", GRF29_4_buffer[clk]);
        end
        if (GRF29_5_buffer[clk] != GRF29_5_buffer[!clk]) begin
          $fwrite(f, "Register (29,5) Value: %h\n", GRF29_5_buffer[clk]);
        end
        if (GRF29_6_buffer[clk] != GRF29_6_buffer[!clk]) begin
          $fwrite(f, "Register (29,6) Value: %h\n", GRF29_6_buffer[clk]);
        end
        if (GRF29_7_buffer[clk] != GRF29_7_buffer[!clk]) begin
          $fwrite(f, "Register (29,7) Value: %h\n", GRF29_7_buffer[clk]);
        end
        if (GRF29_8_buffer[clk] != GRF29_8_buffer[!clk]) begin
          $fwrite(f, "Register (29,8) Value: %h\n", GRF29_8_buffer[clk]);
        end
        if (GRF29_9_buffer[clk] != GRF29_9_buffer[!clk]) begin
          $fwrite(f, "Register (29,9) Value: %h\n", GRF29_9_buffer[clk]);
        end
        if (GRF29_10_buffer[clk] != GRF29_10_buffer[!clk]) begin
          $fwrite(f, "Register (29,10) Value: %h\n", GRF29_10_buffer[clk]);
        end
        if (GRF29_11_buffer[clk] != GRF29_11_buffer[!clk]) begin
          $fwrite(f, "Register (29,11) Value: %h\n", GRF29_11_buffer[clk]);
        end
        if (GRF29_12_buffer[clk] != GRF29_12_buffer[!clk]) begin
          $fwrite(f, "Register (29,12) Value: %h\n", GRF29_12_buffer[clk]);
        end
        if (GRF29_13_buffer[clk] != GRF29_13_buffer[!clk]) begin
          $fwrite(f, "Register (29,13) Value: %h\n", GRF29_13_buffer[clk]);
        end
        if (GRF29_14_buffer[clk] != GRF29_14_buffer[!clk]) begin
          $fwrite(f, "Register (29,14) Value: %h\n", GRF29_14_buffer[clk]);
        end
        if (GRF29_15_buffer[clk] != GRF29_15_buffer[!clk]) begin
          $fwrite(f, "Register (29,15) Value: %h\n", GRF29_15_buffer[clk]);
        end
        if (GRF29_16_buffer[clk] != GRF29_16_buffer[!clk]) begin
          $fwrite(f, "Register (29,16) Value: %h\n", GRF29_16_buffer[clk]);
        end
        if (GRF29_17_buffer[clk] != GRF29_17_buffer[!clk]) begin
          $fwrite(f, "Register (29,17) Value: %h\n", GRF29_17_buffer[clk]);
        end
        if (GRF29_18_buffer[clk] != GRF29_18_buffer[!clk]) begin
          $fwrite(f, "Register (29,18) Value: %h\n", GRF29_18_buffer[clk]);
        end
        if (GRF29_19_buffer[clk] != GRF29_19_buffer[!clk]) begin
          $fwrite(f, "Register (29,19) Value: %h\n", GRF29_19_buffer[clk]);
        end
        if (GRF29_20_buffer[clk] != GRF29_20_buffer[!clk]) begin
          $fwrite(f, "Register (29,20) Value: %h\n", GRF29_20_buffer[clk]);
        end
        if (GRF29_21_buffer[clk] != GRF29_21_buffer[!clk]) begin
          $fwrite(f, "Register (29,21) Value: %h\n", GRF29_21_buffer[clk]);
        end
        if (GRF29_22_buffer[clk] != GRF29_22_buffer[!clk]) begin
          $fwrite(f, "Register (29,22) Value: %h\n", GRF29_22_buffer[clk]);
        end
        if (GRF29_23_buffer[clk] != GRF29_23_buffer[!clk]) begin
          $fwrite(f, "Register (29,23) Value: %h\n", GRF29_23_buffer[clk]);
        end
        if (GRF29_24_buffer[clk] != GRF29_24_buffer[!clk]) begin
          $fwrite(f, "Register (29,24) Value: %h\n", GRF29_24_buffer[clk]);
        end
        if (GRF29_25_buffer[clk] != GRF29_25_buffer[!clk]) begin
          $fwrite(f, "Register (29,25) Value: %h\n", GRF29_25_buffer[clk]);
        end
        if (GRF29_26_buffer[clk] != GRF29_26_buffer[!clk]) begin
          $fwrite(f, "Register (29,26) Value: %h\n", GRF29_26_buffer[clk]);
        end
        if (GRF29_27_buffer[clk] != GRF29_27_buffer[!clk]) begin
          $fwrite(f, "Register (29,27) Value: %h\n", GRF29_27_buffer[clk]);
        end
        if (GRF29_28_buffer[clk] != GRF29_28_buffer[!clk]) begin
          $fwrite(f, "Register (29,28) Value: %h\n", GRF29_28_buffer[clk]);
        end
        if (GRF29_29_buffer[clk] != GRF29_29_buffer[!clk]) begin
          $fwrite(f, "Register (29,29) Value: %h\n", GRF29_29_buffer[clk]);
        end
        if (GRF29_30_buffer[clk] != GRF29_30_buffer[!clk]) begin
          $fwrite(f, "Register (29,30) Value: %h\n", GRF29_30_buffer[clk]);
        end
        if (GRF29_31_buffer[clk] != GRF29_31_buffer[!clk]) begin
          $fwrite(f, "Register (29,31) Value: %h\n", GRF29_31_buffer[clk]);
        end
        if (GRF30_0_buffer[clk] != GRF30_0_buffer[!clk]) begin
          $fwrite(f, "Register (30,0) Value: %h\n", GRF30_0_buffer[clk]);
        end
        if (GRF30_1_buffer[clk] != GRF30_1_buffer[!clk]) begin
          $fwrite(f, "Register (30,1) Value: %h\n", GRF30_1_buffer[clk]);
        end
        if (GRF30_2_buffer[clk] != GRF30_2_buffer[!clk]) begin
          $fwrite(f, "Register (30,2) Value: %h\n", GRF30_2_buffer[clk]);
        end
        if (GRF30_3_buffer[clk] != GRF30_3_buffer[!clk]) begin
          $fwrite(f, "Register (30,3) Value: %h\n", GRF30_3_buffer[clk]);
        end
        if (GRF30_4_buffer[clk] != GRF30_4_buffer[!clk]) begin
          $fwrite(f, "Register (30,4) Value: %h\n", GRF30_4_buffer[clk]);
        end
        if (GRF30_5_buffer[clk] != GRF30_5_buffer[!clk]) begin
          $fwrite(f, "Register (30,5) Value: %h\n", GRF30_5_buffer[clk]);
        end
        if (GRF30_6_buffer[clk] != GRF30_6_buffer[!clk]) begin
          $fwrite(f, "Register (30,6) Value: %h\n", GRF30_6_buffer[clk]);
        end
        if (GRF30_7_buffer[clk] != GRF30_7_buffer[!clk]) begin
          $fwrite(f, "Register (30,7) Value: %h\n", GRF30_7_buffer[clk]);
        end
        if (GRF30_8_buffer[clk] != GRF30_8_buffer[!clk]) begin
          $fwrite(f, "Register (30,8) Value: %h\n", GRF30_8_buffer[clk]);
        end
        if (GRF30_9_buffer[clk] != GRF30_9_buffer[!clk]) begin
          $fwrite(f, "Register (30,9) Value: %h\n", GRF30_9_buffer[clk]);
        end
        if (GRF30_10_buffer[clk] != GRF30_10_buffer[!clk]) begin
          $fwrite(f, "Register (30,10) Value: %h\n", GRF30_10_buffer[clk]);
        end
        if (GRF30_11_buffer[clk] != GRF30_11_buffer[!clk]) begin
          $fwrite(f, "Register (30,11) Value: %h\n", GRF30_11_buffer[clk]);
        end
        if (GRF30_12_buffer[clk] != GRF30_12_buffer[!clk]) begin
          $fwrite(f, "Register (30,12) Value: %h\n", GRF30_12_buffer[clk]);
        end
        if (GRF30_13_buffer[clk] != GRF30_13_buffer[!clk]) begin
          $fwrite(f, "Register (30,13) Value: %h\n", GRF30_13_buffer[clk]);
        end
        if (GRF30_14_buffer[clk] != GRF30_14_buffer[!clk]) begin
          $fwrite(f, "Register (30,14) Value: %h\n", GRF30_14_buffer[clk]);
        end
        if (GRF30_15_buffer[clk] != GRF30_15_buffer[!clk]) begin
          $fwrite(f, "Register (30,15) Value: %h\n", GRF30_15_buffer[clk]);
        end
        if (GRF30_16_buffer[clk] != GRF30_16_buffer[!clk]) begin
          $fwrite(f, "Register (30,16) Value: %h\n", GRF30_16_buffer[clk]);
        end
        if (GRF30_17_buffer[clk] != GRF30_17_buffer[!clk]) begin
          $fwrite(f, "Register (30,17) Value: %h\n", GRF30_17_buffer[clk]);
        end
        if (GRF30_18_buffer[clk] != GRF30_18_buffer[!clk]) begin
          $fwrite(f, "Register (30,18) Value: %h\n", GRF30_18_buffer[clk]);
        end
        if (GRF30_19_buffer[clk] != GRF30_19_buffer[!clk]) begin
          $fwrite(f, "Register (30,19) Value: %h\n", GRF30_19_buffer[clk]);
        end
        if (GRF30_20_buffer[clk] != GRF30_20_buffer[!clk]) begin
          $fwrite(f, "Register (30,20) Value: %h\n", GRF30_20_buffer[clk]);
        end
        if (GRF30_21_buffer[clk] != GRF30_21_buffer[!clk]) begin
          $fwrite(f, "Register (30,21) Value: %h\n", GRF30_21_buffer[clk]);
        end
        if (GRF30_22_buffer[clk] != GRF30_22_buffer[!clk]) begin
          $fwrite(f, "Register (30,22) Value: %h\n", GRF30_22_buffer[clk]);
        end
        if (GRF30_23_buffer[clk] != GRF30_23_buffer[!clk]) begin
          $fwrite(f, "Register (30,23) Value: %h\n", GRF30_23_buffer[clk]);
        end
        if (GRF30_24_buffer[clk] != GRF30_24_buffer[!clk]) begin
          $fwrite(f, "Register (30,24) Value: %h\n", GRF30_24_buffer[clk]);
        end
        if (GRF30_25_buffer[clk] != GRF30_25_buffer[!clk]) begin
          $fwrite(f, "Register (30,25) Value: %h\n", GRF30_25_buffer[clk]);
        end
        if (GRF30_26_buffer[clk] != GRF30_26_buffer[!clk]) begin
          $fwrite(f, "Register (30,26) Value: %h\n", GRF30_26_buffer[clk]);
        end
        if (GRF30_27_buffer[clk] != GRF30_27_buffer[!clk]) begin
          $fwrite(f, "Register (30,27) Value: %h\n", GRF30_27_buffer[clk]);
        end
        if (GRF30_28_buffer[clk] != GRF30_28_buffer[!clk]) begin
          $fwrite(f, "Register (30,28) Value: %h\n", GRF30_28_buffer[clk]);
        end
        if (GRF30_29_buffer[clk] != GRF30_29_buffer[!clk]) begin
          $fwrite(f, "Register (30,29) Value: %h\n", GRF30_29_buffer[clk]);
        end
        if (GRF30_30_buffer[clk] != GRF30_30_buffer[!clk]) begin
          $fwrite(f, "Register (30,30) Value: %h\n", GRF30_30_buffer[clk]);
        end
        if (GRF30_31_buffer[clk] != GRF30_31_buffer[!clk]) begin
          $fwrite(f, "Register (30,31) Value: %h\n", GRF30_31_buffer[clk]);
        end
        if (GRF31_0_buffer[clk] != GRF31_0_buffer[!clk]) begin
          $fwrite(f, "Register (31,0) Value: %h\n", GRF31_0_buffer[clk]);
        end
        if (GRF31_1_buffer[clk] != GRF31_1_buffer[!clk]) begin
          $fwrite(f, "Register (31,1) Value: %h\n", GRF31_1_buffer[clk]);
        end
        if (GRF31_2_buffer[clk] != GRF31_2_buffer[!clk]) begin
          $fwrite(f, "Register (31,2) Value: %h\n", GRF31_2_buffer[clk]);
        end
        if (GRF31_3_buffer[clk] != GRF31_3_buffer[!clk]) begin
          $fwrite(f, "Register (31,3) Value: %h\n", GRF31_3_buffer[clk]);
        end
        if (GRF31_4_buffer[clk] != GRF31_4_buffer[!clk]) begin
          $fwrite(f, "Register (31,4) Value: %h\n", GRF31_4_buffer[clk]);
        end
        if (GRF31_5_buffer[clk] != GRF31_5_buffer[!clk]) begin
          $fwrite(f, "Register (31,5) Value: %h\n", GRF31_5_buffer[clk]);
        end
        if (GRF31_6_buffer[clk] != GRF31_6_buffer[!clk]) begin
          $fwrite(f, "Register (31,6) Value: %h\n", GRF31_6_buffer[clk]);
        end
        if (GRF31_7_buffer[clk] != GRF31_7_buffer[!clk]) begin
          $fwrite(f, "Register (31,7) Value: %h\n", GRF31_7_buffer[clk]);
        end
        if (GRF31_8_buffer[clk] != GRF31_8_buffer[!clk]) begin
          $fwrite(f, "Register (31,8) Value: %h\n", GRF31_8_buffer[clk]);
        end
        if (GRF31_9_buffer[clk] != GRF31_9_buffer[!clk]) begin
          $fwrite(f, "Register (31,9) Value: %h\n", GRF31_9_buffer[clk]);
        end
        if (GRF31_10_buffer[clk] != GRF31_10_buffer[!clk]) begin
          $fwrite(f, "Register (31,10) Value: %h\n", GRF31_10_buffer[clk]);
        end
        if (GRF31_11_buffer[clk] != GRF31_11_buffer[!clk]) begin
          $fwrite(f, "Register (31,11) Value: %h\n", GRF31_11_buffer[clk]);
        end
        if (GRF31_12_buffer[clk] != GRF31_12_buffer[!clk]) begin
          $fwrite(f, "Register (31,12) Value: %h\n", GRF31_12_buffer[clk]);
        end
        if (GRF31_13_buffer[clk] != GRF31_13_buffer[!clk]) begin
          $fwrite(f, "Register (31,13) Value: %h\n", GRF31_13_buffer[clk]);
        end
        if (GRF31_14_buffer[clk] != GRF31_14_buffer[!clk]) begin
          $fwrite(f, "Register (31,14) Value: %h\n", GRF31_14_buffer[clk]);
        end
        if (GRF31_15_buffer[clk] != GRF31_15_buffer[!clk]) begin
          $fwrite(f, "Register (31,15) Value: %h\n", GRF31_15_buffer[clk]);
        end
        if (GRF31_16_buffer[clk] != GRF31_16_buffer[!clk]) begin
          $fwrite(f, "Register (31,16) Value: %h\n", GRF31_16_buffer[clk]);
        end
        if (GRF31_17_buffer[clk] != GRF31_17_buffer[!clk]) begin
          $fwrite(f, "Register (31,17) Value: %h\n", GRF31_17_buffer[clk]);
        end
        if (GRF31_18_buffer[clk] != GRF31_18_buffer[!clk]) begin
          $fwrite(f, "Register (31,18) Value: %h\n", GRF31_18_buffer[clk]);
        end
        if (GRF31_19_buffer[clk] != GRF31_19_buffer[!clk]) begin
          $fwrite(f, "Register (31,19) Value: %h\n", GRF31_19_buffer[clk]);
        end
        if (GRF31_20_buffer[clk] != GRF31_20_buffer[!clk]) begin
          $fwrite(f, "Register (31,20) Value: %h\n", GRF31_20_buffer[clk]);
        end
        if (GRF31_21_buffer[clk] != GRF31_21_buffer[!clk]) begin
          $fwrite(f, "Register (31,21) Value: %h\n", GRF31_21_buffer[clk]);
        end
        if (GRF31_22_buffer[clk] != GRF31_22_buffer[!clk]) begin
          $fwrite(f, "Register (31,22) Value: %h\n", GRF31_22_buffer[clk]);
        end
        if (GRF31_23_buffer[clk] != GRF31_23_buffer[!clk]) begin
          $fwrite(f, "Register (31,23) Value: %h\n", GRF31_23_buffer[clk]);
        end
        if (GRF31_24_buffer[clk] != GRF31_24_buffer[!clk]) begin
          $fwrite(f, "Register (31,24) Value: %h\n", GRF31_24_buffer[clk]);
        end
        if (GRF31_25_buffer[clk] != GRF31_25_buffer[!clk]) begin
          $fwrite(f, "Register (31,25) Value: %h\n", GRF31_25_buffer[clk]);
        end
        if (GRF31_26_buffer[clk] != GRF31_26_buffer[!clk]) begin
          $fwrite(f, "Register (31,26) Value: %h\n", GRF31_26_buffer[clk]);
        end
        if (GRF31_27_buffer[clk] != GRF31_27_buffer[!clk]) begin
          $fwrite(f, "Register (31,27) Value: %h\n", GRF31_27_buffer[clk]);
        end
        if (GRF31_28_buffer[clk] != GRF31_28_buffer[!clk]) begin
          $fwrite(f, "Register (31,28) Value: %h\n", GRF31_28_buffer[clk]);
        end
        if (GRF31_29_buffer[clk] != GRF31_29_buffer[!clk]) begin
          $fwrite(f, "Register (31,29) Value: %h\n", GRF31_29_buffer[clk]);
        end
        if (GRF31_30_buffer[clk] != GRF31_30_buffer[!clk]) begin
          $fwrite(f, "Register (31,30) Value: %h\n", GRF31_30_buffer[clk]);
        end
        if (GRF31_31_buffer[clk] != GRF31_31_buffer[!clk]) begin
          $fwrite(f, "Register (31,31) Value: %h\n", GRF31_31_buffer[clk]);
        end
        if (GRF32_0_buffer[clk] != GRF32_0_buffer[!clk]) begin
          $fwrite(f, "Register (32,0) Value: %h\n", GRF32_0_buffer[clk]);
        end
        if (GRF32_1_buffer[clk] != GRF32_1_buffer[!clk]) begin
          $fwrite(f, "Register (32,1) Value: %h\n", GRF32_1_buffer[clk]);
        end
        if (GRF32_2_buffer[clk] != GRF32_2_buffer[!clk]) begin
          $fwrite(f, "Register (32,2) Value: %h\n", GRF32_2_buffer[clk]);
        end
        if (GRF32_3_buffer[clk] != GRF32_3_buffer[!clk]) begin
          $fwrite(f, "Register (32,3) Value: %h\n", GRF32_3_buffer[clk]);
        end
        if (GRF32_4_buffer[clk] != GRF32_4_buffer[!clk]) begin
          $fwrite(f, "Register (32,4) Value: %h\n", GRF32_4_buffer[clk]);
        end
        if (GRF32_5_buffer[clk] != GRF32_5_buffer[!clk]) begin
          $fwrite(f, "Register (32,5) Value: %h\n", GRF32_5_buffer[clk]);
        end
        if (GRF32_6_buffer[clk] != GRF32_6_buffer[!clk]) begin
          $fwrite(f, "Register (32,6) Value: %h\n", GRF32_6_buffer[clk]);
        end
        if (GRF32_7_buffer[clk] != GRF32_7_buffer[!clk]) begin
          $fwrite(f, "Register (32,7) Value: %h\n", GRF32_7_buffer[clk]);
        end
        if (GRF32_8_buffer[clk] != GRF32_8_buffer[!clk]) begin
          $fwrite(f, "Register (32,8) Value: %h\n", GRF32_8_buffer[clk]);
        end
        if (GRF32_9_buffer[clk] != GRF32_9_buffer[!clk]) begin
          $fwrite(f, "Register (32,9) Value: %h\n", GRF32_9_buffer[clk]);
        end
        if (GRF32_10_buffer[clk] != GRF32_10_buffer[!clk]) begin
          $fwrite(f, "Register (32,10) Value: %h\n", GRF32_10_buffer[clk]);
        end
        if (GRF32_11_buffer[clk] != GRF32_11_buffer[!clk]) begin
          $fwrite(f, "Register (32,11) Value: %h\n", GRF32_11_buffer[clk]);
        end
        if (GRF32_12_buffer[clk] != GRF32_12_buffer[!clk]) begin
          $fwrite(f, "Register (32,12) Value: %h\n", GRF32_12_buffer[clk]);
        end
        if (GRF32_13_buffer[clk] != GRF32_13_buffer[!clk]) begin
          $fwrite(f, "Register (32,13) Value: %h\n", GRF32_13_buffer[clk]);
        end
        if (GRF32_14_buffer[clk] != GRF32_14_buffer[!clk]) begin
          $fwrite(f, "Register (32,14) Value: %h\n", GRF32_14_buffer[clk]);
        end
        if (GRF32_15_buffer[clk] != GRF32_15_buffer[!clk]) begin
          $fwrite(f, "Register (32,15) Value: %h\n", GRF32_15_buffer[clk]);
        end
        if (GRF32_16_buffer[clk] != GRF32_16_buffer[!clk]) begin
          $fwrite(f, "Register (32,16) Value: %h\n", GRF32_16_buffer[clk]);
        end
        if (GRF32_17_buffer[clk] != GRF32_17_buffer[!clk]) begin
          $fwrite(f, "Register (32,17) Value: %h\n", GRF32_17_buffer[clk]);
        end
        if (GRF32_18_buffer[clk] != GRF32_18_buffer[!clk]) begin
          $fwrite(f, "Register (32,18) Value: %h\n", GRF32_18_buffer[clk]);
        end
        if (GRF32_19_buffer[clk] != GRF32_19_buffer[!clk]) begin
          $fwrite(f, "Register (32,19) Value: %h\n", GRF32_19_buffer[clk]);
        end
        if (GRF32_20_buffer[clk] != GRF32_20_buffer[!clk]) begin
          $fwrite(f, "Register (32,20) Value: %h\n", GRF32_20_buffer[clk]);
        end
        if (GRF32_21_buffer[clk] != GRF32_21_buffer[!clk]) begin
          $fwrite(f, "Register (32,21) Value: %h\n", GRF32_21_buffer[clk]);
        end
        if (GRF32_22_buffer[clk] != GRF32_22_buffer[!clk]) begin
          $fwrite(f, "Register (32,22) Value: %h\n", GRF32_22_buffer[clk]);
        end
        if (GRF32_23_buffer[clk] != GRF32_23_buffer[!clk]) begin
          $fwrite(f, "Register (32,23) Value: %h\n", GRF32_23_buffer[clk]);
        end
        if (GRF32_24_buffer[clk] != GRF32_24_buffer[!clk]) begin
          $fwrite(f, "Register (32,24) Value: %h\n", GRF32_24_buffer[clk]);
        end
        if (GRF32_25_buffer[clk] != GRF32_25_buffer[!clk]) begin
          $fwrite(f, "Register (32,25) Value: %h\n", GRF32_25_buffer[clk]);
        end
        if (GRF32_26_buffer[clk] != GRF32_26_buffer[!clk]) begin
          $fwrite(f, "Register (32,26) Value: %h\n", GRF32_26_buffer[clk]);
        end
        if (GRF32_27_buffer[clk] != GRF32_27_buffer[!clk]) begin
          $fwrite(f, "Register (32,27) Value: %h\n", GRF32_27_buffer[clk]);
        end
        if (GRF32_28_buffer[clk] != GRF32_28_buffer[!clk]) begin
          $fwrite(f, "Register (32,28) Value: %h\n", GRF32_28_buffer[clk]);
        end
        if (GRF32_29_buffer[clk] != GRF32_29_buffer[!clk]) begin
          $fwrite(f, "Register (32,29) Value: %h\n", GRF32_29_buffer[clk]);
        end
        if (GRF32_30_buffer[clk] != GRF32_30_buffer[!clk]) begin
          $fwrite(f, "Register (32,30) Value: %h\n", GRF32_30_buffer[clk]);
        end
        if (GRF32_31_buffer[clk] != GRF32_31_buffer[!clk]) begin
          $fwrite(f, "Register (32,31) Value: %h\n", GRF32_31_buffer[clk]);
        end
        if (GRF33_0_buffer[clk] != GRF33_0_buffer[!clk]) begin
          $fwrite(f, "Register (33,0) Value: %h\n", GRF33_0_buffer[clk]);
        end
        if (GRF33_1_buffer[clk] != GRF33_1_buffer[!clk]) begin
          $fwrite(f, "Register (33,1) Value: %h\n", GRF33_1_buffer[clk]);
        end
        if (GRF33_2_buffer[clk] != GRF33_2_buffer[!clk]) begin
          $fwrite(f, "Register (33,2) Value: %h\n", GRF33_2_buffer[clk]);
        end
        if (GRF33_3_buffer[clk] != GRF33_3_buffer[!clk]) begin
          $fwrite(f, "Register (33,3) Value: %h\n", GRF33_3_buffer[clk]);
        end
        if (GRF33_4_buffer[clk] != GRF33_4_buffer[!clk]) begin
          $fwrite(f, "Register (33,4) Value: %h\n", GRF33_4_buffer[clk]);
        end
        if (GRF33_5_buffer[clk] != GRF33_5_buffer[!clk]) begin
          $fwrite(f, "Register (33,5) Value: %h\n", GRF33_5_buffer[clk]);
        end
        if (GRF33_6_buffer[clk] != GRF33_6_buffer[!clk]) begin
          $fwrite(f, "Register (33,6) Value: %h\n", GRF33_6_buffer[clk]);
        end
        if (GRF33_7_buffer[clk] != GRF33_7_buffer[!clk]) begin
          $fwrite(f, "Register (33,7) Value: %h\n", GRF33_7_buffer[clk]);
        end
        if (GRF33_8_buffer[clk] != GRF33_8_buffer[!clk]) begin
          $fwrite(f, "Register (33,8) Value: %h\n", GRF33_8_buffer[clk]);
        end
        if (GRF33_9_buffer[clk] != GRF33_9_buffer[!clk]) begin
          $fwrite(f, "Register (33,9) Value: %h\n", GRF33_9_buffer[clk]);
        end
        if (GRF33_10_buffer[clk] != GRF33_10_buffer[!clk]) begin
          $fwrite(f, "Register (33,10) Value: %h\n", GRF33_10_buffer[clk]);
        end
        if (GRF33_11_buffer[clk] != GRF33_11_buffer[!clk]) begin
          $fwrite(f, "Register (33,11) Value: %h\n", GRF33_11_buffer[clk]);
        end
        if (GRF33_12_buffer[clk] != GRF33_12_buffer[!clk]) begin
          $fwrite(f, "Register (33,12) Value: %h\n", GRF33_12_buffer[clk]);
        end
        if (GRF33_13_buffer[clk] != GRF33_13_buffer[!clk]) begin
          $fwrite(f, "Register (33,13) Value: %h\n", GRF33_13_buffer[clk]);
        end
        if (GRF33_14_buffer[clk] != GRF33_14_buffer[!clk]) begin
          $fwrite(f, "Register (33,14) Value: %h\n", GRF33_14_buffer[clk]);
        end
        if (GRF33_15_buffer[clk] != GRF33_15_buffer[!clk]) begin
          $fwrite(f, "Register (33,15) Value: %h\n", GRF33_15_buffer[clk]);
        end
        if (GRF33_16_buffer[clk] != GRF33_16_buffer[!clk]) begin
          $fwrite(f, "Register (33,16) Value: %h\n", GRF33_16_buffer[clk]);
        end
        if (GRF33_17_buffer[clk] != GRF33_17_buffer[!clk]) begin
          $fwrite(f, "Register (33,17) Value: %h\n", GRF33_17_buffer[clk]);
        end
        if (GRF33_18_buffer[clk] != GRF33_18_buffer[!clk]) begin
          $fwrite(f, "Register (33,18) Value: %h\n", GRF33_18_buffer[clk]);
        end
        if (GRF33_19_buffer[clk] != GRF33_19_buffer[!clk]) begin
          $fwrite(f, "Register (33,19) Value: %h\n", GRF33_19_buffer[clk]);
        end
        if (GRF33_20_buffer[clk] != GRF33_20_buffer[!clk]) begin
          $fwrite(f, "Register (33,20) Value: %h\n", GRF33_20_buffer[clk]);
        end
        if (GRF33_21_buffer[clk] != GRF33_21_buffer[!clk]) begin
          $fwrite(f, "Register (33,21) Value: %h\n", GRF33_21_buffer[clk]);
        end
        if (GRF33_22_buffer[clk] != GRF33_22_buffer[!clk]) begin
          $fwrite(f, "Register (33,22) Value: %h\n", GRF33_22_buffer[clk]);
        end
        if (GRF33_23_buffer[clk] != GRF33_23_buffer[!clk]) begin
          $fwrite(f, "Register (33,23) Value: %h\n", GRF33_23_buffer[clk]);
        end
        if (GRF33_24_buffer[clk] != GRF33_24_buffer[!clk]) begin
          $fwrite(f, "Register (33,24) Value: %h\n", GRF33_24_buffer[clk]);
        end
        if (GRF33_25_buffer[clk] != GRF33_25_buffer[!clk]) begin
          $fwrite(f, "Register (33,25) Value: %h\n", GRF33_25_buffer[clk]);
        end
        if (GRF33_26_buffer[clk] != GRF33_26_buffer[!clk]) begin
          $fwrite(f, "Register (33,26) Value: %h\n", GRF33_26_buffer[clk]);
        end
        if (GRF33_27_buffer[clk] != GRF33_27_buffer[!clk]) begin
          $fwrite(f, "Register (33,27) Value: %h\n", GRF33_27_buffer[clk]);
        end
        if (GRF33_28_buffer[clk] != GRF33_28_buffer[!clk]) begin
          $fwrite(f, "Register (33,28) Value: %h\n", GRF33_28_buffer[clk]);
        end
        if (GRF33_29_buffer[clk] != GRF33_29_buffer[!clk]) begin
          $fwrite(f, "Register (33,29) Value: %h\n", GRF33_29_buffer[clk]);
        end
        if (GRF33_30_buffer[clk] != GRF33_30_buffer[!clk]) begin
          $fwrite(f, "Register (33,30) Value: %h\n", GRF33_30_buffer[clk]);
        end
        if (GRF33_31_buffer[clk] != GRF33_31_buffer[!clk]) begin
          $fwrite(f, "Register (33,31) Value: %h\n", GRF33_31_buffer[clk]);
        end
        if (GRF34_0_buffer[clk] != GRF34_0_buffer[!clk]) begin
          $fwrite(f, "Register (34,0) Value: %h\n", GRF34_0_buffer[clk]);
        end
        if (GRF34_1_buffer[clk] != GRF34_1_buffer[!clk]) begin
          $fwrite(f, "Register (34,1) Value: %h\n", GRF34_1_buffer[clk]);
        end
        if (GRF34_2_buffer[clk] != GRF34_2_buffer[!clk]) begin
          $fwrite(f, "Register (34,2) Value: %h\n", GRF34_2_buffer[clk]);
        end
        if (GRF34_3_buffer[clk] != GRF34_3_buffer[!clk]) begin
          $fwrite(f, "Register (34,3) Value: %h\n", GRF34_3_buffer[clk]);
        end
        if (GRF34_4_buffer[clk] != GRF34_4_buffer[!clk]) begin
          $fwrite(f, "Register (34,4) Value: %h\n", GRF34_4_buffer[clk]);
        end
        if (GRF34_5_buffer[clk] != GRF34_5_buffer[!clk]) begin
          $fwrite(f, "Register (34,5) Value: %h\n", GRF34_5_buffer[clk]);
        end
        if (GRF34_6_buffer[clk] != GRF34_6_buffer[!clk]) begin
          $fwrite(f, "Register (34,6) Value: %h\n", GRF34_6_buffer[clk]);
        end
        if (GRF34_7_buffer[clk] != GRF34_7_buffer[!clk]) begin
          $fwrite(f, "Register (34,7) Value: %h\n", GRF34_7_buffer[clk]);
        end
        if (GRF34_8_buffer[clk] != GRF34_8_buffer[!clk]) begin
          $fwrite(f, "Register (34,8) Value: %h\n", GRF34_8_buffer[clk]);
        end
        if (GRF34_9_buffer[clk] != GRF34_9_buffer[!clk]) begin
          $fwrite(f, "Register (34,9) Value: %h\n", GRF34_9_buffer[clk]);
        end
        if (GRF34_10_buffer[clk] != GRF34_10_buffer[!clk]) begin
          $fwrite(f, "Register (34,10) Value: %h\n", GRF34_10_buffer[clk]);
        end
        if (GRF34_11_buffer[clk] != GRF34_11_buffer[!clk]) begin
          $fwrite(f, "Register (34,11) Value: %h\n", GRF34_11_buffer[clk]);
        end
        if (GRF34_12_buffer[clk] != GRF34_12_buffer[!clk]) begin
          $fwrite(f, "Register (34,12) Value: %h\n", GRF34_12_buffer[clk]);
        end
        if (GRF34_13_buffer[clk] != GRF34_13_buffer[!clk]) begin
          $fwrite(f, "Register (34,13) Value: %h\n", GRF34_13_buffer[clk]);
        end
        if (GRF34_14_buffer[clk] != GRF34_14_buffer[!clk]) begin
          $fwrite(f, "Register (34,14) Value: %h\n", GRF34_14_buffer[clk]);
        end
        if (GRF34_15_buffer[clk] != GRF34_15_buffer[!clk]) begin
          $fwrite(f, "Register (34,15) Value: %h\n", GRF34_15_buffer[clk]);
        end
        if (GRF34_16_buffer[clk] != GRF34_16_buffer[!clk]) begin
          $fwrite(f, "Register (34,16) Value: %h\n", GRF34_16_buffer[clk]);
        end
        if (GRF34_17_buffer[clk] != GRF34_17_buffer[!clk]) begin
          $fwrite(f, "Register (34,17) Value: %h\n", GRF34_17_buffer[clk]);
        end
        if (GRF34_18_buffer[clk] != GRF34_18_buffer[!clk]) begin
          $fwrite(f, "Register (34,18) Value: %h\n", GRF34_18_buffer[clk]);
        end
        if (GRF34_19_buffer[clk] != GRF34_19_buffer[!clk]) begin
          $fwrite(f, "Register (34,19) Value: %h\n", GRF34_19_buffer[clk]);
        end
        if (GRF34_20_buffer[clk] != GRF34_20_buffer[!clk]) begin
          $fwrite(f, "Register (34,20) Value: %h\n", GRF34_20_buffer[clk]);
        end
        if (GRF34_21_buffer[clk] != GRF34_21_buffer[!clk]) begin
          $fwrite(f, "Register (34,21) Value: %h\n", GRF34_21_buffer[clk]);
        end
        if (GRF34_22_buffer[clk] != GRF34_22_buffer[!clk]) begin
          $fwrite(f, "Register (34,22) Value: %h\n", GRF34_22_buffer[clk]);
        end
        if (GRF34_23_buffer[clk] != GRF34_23_buffer[!clk]) begin
          $fwrite(f, "Register (34,23) Value: %h\n", GRF34_23_buffer[clk]);
        end
        if (GRF34_24_buffer[clk] != GRF34_24_buffer[!clk]) begin
          $fwrite(f, "Register (34,24) Value: %h\n", GRF34_24_buffer[clk]);
        end
        if (GRF34_25_buffer[clk] != GRF34_25_buffer[!clk]) begin
          $fwrite(f, "Register (34,25) Value: %h\n", GRF34_25_buffer[clk]);
        end
        if (GRF34_26_buffer[clk] != GRF34_26_buffer[!clk]) begin
          $fwrite(f, "Register (34,26) Value: %h\n", GRF34_26_buffer[clk]);
        end
        if (GRF34_27_buffer[clk] != GRF34_27_buffer[!clk]) begin
          $fwrite(f, "Register (34,27) Value: %h\n", GRF34_27_buffer[clk]);
        end
        if (GRF34_28_buffer[clk] != GRF34_28_buffer[!clk]) begin
          $fwrite(f, "Register (34,28) Value: %h\n", GRF34_28_buffer[clk]);
        end
        if (GRF34_29_buffer[clk] != GRF34_29_buffer[!clk]) begin
          $fwrite(f, "Register (34,29) Value: %h\n", GRF34_29_buffer[clk]);
        end
        if (GRF34_30_buffer[clk] != GRF34_30_buffer[!clk]) begin
          $fwrite(f, "Register (34,30) Value: %h\n", GRF34_30_buffer[clk]);
        end
        if (GRF34_31_buffer[clk] != GRF34_31_buffer[!clk]) begin
          $fwrite(f, "Register (34,31) Value: %h\n", GRF34_31_buffer[clk]);
        end
        if (GRF35_0_buffer[clk] != GRF35_0_buffer[!clk]) begin
          $fwrite(f, "Register (35,0) Value: %h\n", GRF35_0_buffer[clk]);
        end
        if (GRF35_1_buffer[clk] != GRF35_1_buffer[!clk]) begin
          $fwrite(f, "Register (35,1) Value: %h\n", GRF35_1_buffer[clk]);
        end
        if (GRF35_2_buffer[clk] != GRF35_2_buffer[!clk]) begin
          $fwrite(f, "Register (35,2) Value: %h\n", GRF35_2_buffer[clk]);
        end
        if (GRF35_3_buffer[clk] != GRF35_3_buffer[!clk]) begin
          $fwrite(f, "Register (35,3) Value: %h\n", GRF35_3_buffer[clk]);
        end
        if (GRF35_4_buffer[clk] != GRF35_4_buffer[!clk]) begin
          $fwrite(f, "Register (35,4) Value: %h\n", GRF35_4_buffer[clk]);
        end
        if (GRF35_5_buffer[clk] != GRF35_5_buffer[!clk]) begin
          $fwrite(f, "Register (35,5) Value: %h\n", GRF35_5_buffer[clk]);
        end
        if (GRF35_6_buffer[clk] != GRF35_6_buffer[!clk]) begin
          $fwrite(f, "Register (35,6) Value: %h\n", GRF35_6_buffer[clk]);
        end
        if (GRF35_7_buffer[clk] != GRF35_7_buffer[!clk]) begin
          $fwrite(f, "Register (35,7) Value: %h\n", GRF35_7_buffer[clk]);
        end
        if (GRF35_8_buffer[clk] != GRF35_8_buffer[!clk]) begin
          $fwrite(f, "Register (35,8) Value: %h\n", GRF35_8_buffer[clk]);
        end
        if (GRF35_9_buffer[clk] != GRF35_9_buffer[!clk]) begin
          $fwrite(f, "Register (35,9) Value: %h\n", GRF35_9_buffer[clk]);
        end
        if (GRF35_10_buffer[clk] != GRF35_10_buffer[!clk]) begin
          $fwrite(f, "Register (35,10) Value: %h\n", GRF35_10_buffer[clk]);
        end
        if (GRF35_11_buffer[clk] != GRF35_11_buffer[!clk]) begin
          $fwrite(f, "Register (35,11) Value: %h\n", GRF35_11_buffer[clk]);
        end
        if (GRF35_12_buffer[clk] != GRF35_12_buffer[!clk]) begin
          $fwrite(f, "Register (35,12) Value: %h\n", GRF35_12_buffer[clk]);
        end
        if (GRF35_13_buffer[clk] != GRF35_13_buffer[!clk]) begin
          $fwrite(f, "Register (35,13) Value: %h\n", GRF35_13_buffer[clk]);
        end
        if (GRF35_14_buffer[clk] != GRF35_14_buffer[!clk]) begin
          $fwrite(f, "Register (35,14) Value: %h\n", GRF35_14_buffer[clk]);
        end
        if (GRF35_15_buffer[clk] != GRF35_15_buffer[!clk]) begin
          $fwrite(f, "Register (35,15) Value: %h\n", GRF35_15_buffer[clk]);
        end
        if (GRF35_16_buffer[clk] != GRF35_16_buffer[!clk]) begin
          $fwrite(f, "Register (35,16) Value: %h\n", GRF35_16_buffer[clk]);
        end
        if (GRF35_17_buffer[clk] != GRF35_17_buffer[!clk]) begin
          $fwrite(f, "Register (35,17) Value: %h\n", GRF35_17_buffer[clk]);
        end
        if (GRF35_18_buffer[clk] != GRF35_18_buffer[!clk]) begin
          $fwrite(f, "Register (35,18) Value: %h\n", GRF35_18_buffer[clk]);
        end
        if (GRF35_19_buffer[clk] != GRF35_19_buffer[!clk]) begin
          $fwrite(f, "Register (35,19) Value: %h\n", GRF35_19_buffer[clk]);
        end
        if (GRF35_20_buffer[clk] != GRF35_20_buffer[!clk]) begin
          $fwrite(f, "Register (35,20) Value: %h\n", GRF35_20_buffer[clk]);
        end
        if (GRF35_21_buffer[clk] != GRF35_21_buffer[!clk]) begin
          $fwrite(f, "Register (35,21) Value: %h\n", GRF35_21_buffer[clk]);
        end
        if (GRF35_22_buffer[clk] != GRF35_22_buffer[!clk]) begin
          $fwrite(f, "Register (35,22) Value: %h\n", GRF35_22_buffer[clk]);
        end
        if (GRF35_23_buffer[clk] != GRF35_23_buffer[!clk]) begin
          $fwrite(f, "Register (35,23) Value: %h\n", GRF35_23_buffer[clk]);
        end
        if (GRF35_24_buffer[clk] != GRF35_24_buffer[!clk]) begin
          $fwrite(f, "Register (35,24) Value: %h\n", GRF35_24_buffer[clk]);
        end
        if (GRF35_25_buffer[clk] != GRF35_25_buffer[!clk]) begin
          $fwrite(f, "Register (35,25) Value: %h\n", GRF35_25_buffer[clk]);
        end
        if (GRF35_26_buffer[clk] != GRF35_26_buffer[!clk]) begin
          $fwrite(f, "Register (35,26) Value: %h\n", GRF35_26_buffer[clk]);
        end
        if (GRF35_27_buffer[clk] != GRF35_27_buffer[!clk]) begin
          $fwrite(f, "Register (35,27) Value: %h\n", GRF35_27_buffer[clk]);
        end
        if (GRF35_28_buffer[clk] != GRF35_28_buffer[!clk]) begin
          $fwrite(f, "Register (35,28) Value: %h\n", GRF35_28_buffer[clk]);
        end
        if (GRF35_29_buffer[clk] != GRF35_29_buffer[!clk]) begin
          $fwrite(f, "Register (35,29) Value: %h\n", GRF35_29_buffer[clk]);
        end
        if (GRF35_30_buffer[clk] != GRF35_30_buffer[!clk]) begin
          $fwrite(f, "Register (35,30) Value: %h\n", GRF35_30_buffer[clk]);
        end
        if (GRF35_31_buffer[clk] != GRF35_31_buffer[!clk]) begin
          $fwrite(f, "Register (35,31) Value: %h\n", GRF35_31_buffer[clk]);
        end
        if (GRF36_0_buffer[clk] != GRF36_0_buffer[!clk]) begin
          $fwrite(f, "Register (36,0) Value: %h\n", GRF36_0_buffer[clk]);
        end
        if (GRF36_1_buffer[clk] != GRF36_1_buffer[!clk]) begin
          $fwrite(f, "Register (36,1) Value: %h\n", GRF36_1_buffer[clk]);
        end
        if (GRF36_2_buffer[clk] != GRF36_2_buffer[!clk]) begin
          $fwrite(f, "Register (36,2) Value: %h\n", GRF36_2_buffer[clk]);
        end
        if (GRF36_3_buffer[clk] != GRF36_3_buffer[!clk]) begin
          $fwrite(f, "Register (36,3) Value: %h\n", GRF36_3_buffer[clk]);
        end
        if (GRF36_4_buffer[clk] != GRF36_4_buffer[!clk]) begin
          $fwrite(f, "Register (36,4) Value: %h\n", GRF36_4_buffer[clk]);
        end
        if (GRF36_5_buffer[clk] != GRF36_5_buffer[!clk]) begin
          $fwrite(f, "Register (36,5) Value: %h\n", GRF36_5_buffer[clk]);
        end
        if (GRF36_6_buffer[clk] != GRF36_6_buffer[!clk]) begin
          $fwrite(f, "Register (36,6) Value: %h\n", GRF36_6_buffer[clk]);
        end
        if (GRF36_7_buffer[clk] != GRF36_7_buffer[!clk]) begin
          $fwrite(f, "Register (36,7) Value: %h\n", GRF36_7_buffer[clk]);
        end
        if (GRF36_8_buffer[clk] != GRF36_8_buffer[!clk]) begin
          $fwrite(f, "Register (36,8) Value: %h\n", GRF36_8_buffer[clk]);
        end
        if (GRF36_9_buffer[clk] != GRF36_9_buffer[!clk]) begin
          $fwrite(f, "Register (36,9) Value: %h\n", GRF36_9_buffer[clk]);
        end
        if (GRF36_10_buffer[clk] != GRF36_10_buffer[!clk]) begin
          $fwrite(f, "Register (36,10) Value: %h\n", GRF36_10_buffer[clk]);
        end
        if (GRF36_11_buffer[clk] != GRF36_11_buffer[!clk]) begin
          $fwrite(f, "Register (36,11) Value: %h\n", GRF36_11_buffer[clk]);
        end
        if (GRF36_12_buffer[clk] != GRF36_12_buffer[!clk]) begin
          $fwrite(f, "Register (36,12) Value: %h\n", GRF36_12_buffer[clk]);
        end
        if (GRF36_13_buffer[clk] != GRF36_13_buffer[!clk]) begin
          $fwrite(f, "Register (36,13) Value: %h\n", GRF36_13_buffer[clk]);
        end
        if (GRF36_14_buffer[clk] != GRF36_14_buffer[!clk]) begin
          $fwrite(f, "Register (36,14) Value: %h\n", GRF36_14_buffer[clk]);
        end
        if (GRF36_15_buffer[clk] != GRF36_15_buffer[!clk]) begin
          $fwrite(f, "Register (36,15) Value: %h\n", GRF36_15_buffer[clk]);
        end
        if (GRF36_16_buffer[clk] != GRF36_16_buffer[!clk]) begin
          $fwrite(f, "Register (36,16) Value: %h\n", GRF36_16_buffer[clk]);
        end
        if (GRF36_17_buffer[clk] != GRF36_17_buffer[!clk]) begin
          $fwrite(f, "Register (36,17) Value: %h\n", GRF36_17_buffer[clk]);
        end
        if (GRF36_18_buffer[clk] != GRF36_18_buffer[!clk]) begin
          $fwrite(f, "Register (36,18) Value: %h\n", GRF36_18_buffer[clk]);
        end
        if (GRF36_19_buffer[clk] != GRF36_19_buffer[!clk]) begin
          $fwrite(f, "Register (36,19) Value: %h\n", GRF36_19_buffer[clk]);
        end
        if (GRF36_20_buffer[clk] != GRF36_20_buffer[!clk]) begin
          $fwrite(f, "Register (36,20) Value: %h\n", GRF36_20_buffer[clk]);
        end
        if (GRF36_21_buffer[clk] != GRF36_21_buffer[!clk]) begin
          $fwrite(f, "Register (36,21) Value: %h\n", GRF36_21_buffer[clk]);
        end
        if (GRF36_22_buffer[clk] != GRF36_22_buffer[!clk]) begin
          $fwrite(f, "Register (36,22) Value: %h\n", GRF36_22_buffer[clk]);
        end
        if (GRF36_23_buffer[clk] != GRF36_23_buffer[!clk]) begin
          $fwrite(f, "Register (36,23) Value: %h\n", GRF36_23_buffer[clk]);
        end
        if (GRF36_24_buffer[clk] != GRF36_24_buffer[!clk]) begin
          $fwrite(f, "Register (36,24) Value: %h\n", GRF36_24_buffer[clk]);
        end
        if (GRF36_25_buffer[clk] != GRF36_25_buffer[!clk]) begin
          $fwrite(f, "Register (36,25) Value: %h\n", GRF36_25_buffer[clk]);
        end
        if (GRF36_26_buffer[clk] != GRF36_26_buffer[!clk]) begin
          $fwrite(f, "Register (36,26) Value: %h\n", GRF36_26_buffer[clk]);
        end
        if (GRF36_27_buffer[clk] != GRF36_27_buffer[!clk]) begin
          $fwrite(f, "Register (36,27) Value: %h\n", GRF36_27_buffer[clk]);
        end
        if (GRF36_28_buffer[clk] != GRF36_28_buffer[!clk]) begin
          $fwrite(f, "Register (36,28) Value: %h\n", GRF36_28_buffer[clk]);
        end
        if (GRF36_29_buffer[clk] != GRF36_29_buffer[!clk]) begin
          $fwrite(f, "Register (36,29) Value: %h\n", GRF36_29_buffer[clk]);
        end
        if (GRF36_30_buffer[clk] != GRF36_30_buffer[!clk]) begin
          $fwrite(f, "Register (36,30) Value: %h\n", GRF36_30_buffer[clk]);
        end
        if (GRF36_31_buffer[clk] != GRF36_31_buffer[!clk]) begin
          $fwrite(f, "Register (36,31) Value: %h\n", GRF36_31_buffer[clk]);
        end
        if (GRF37_0_buffer[clk] != GRF37_0_buffer[!clk]) begin
          $fwrite(f, "Register (37,0) Value: %h\n", GRF37_0_buffer[clk]);
        end
        if (GRF37_1_buffer[clk] != GRF37_1_buffer[!clk]) begin
          $fwrite(f, "Register (37,1) Value: %h\n", GRF37_1_buffer[clk]);
        end
        if (GRF37_2_buffer[clk] != GRF37_2_buffer[!clk]) begin
          $fwrite(f, "Register (37,2) Value: %h\n", GRF37_2_buffer[clk]);
        end
        if (GRF37_3_buffer[clk] != GRF37_3_buffer[!clk]) begin
          $fwrite(f, "Register (37,3) Value: %h\n", GRF37_3_buffer[clk]);
        end
        if (GRF37_4_buffer[clk] != GRF37_4_buffer[!clk]) begin
          $fwrite(f, "Register (37,4) Value: %h\n", GRF37_4_buffer[clk]);
        end
        if (GRF37_5_buffer[clk] != GRF37_5_buffer[!clk]) begin
          $fwrite(f, "Register (37,5) Value: %h\n", GRF37_5_buffer[clk]);
        end
        if (GRF37_6_buffer[clk] != GRF37_6_buffer[!clk]) begin
          $fwrite(f, "Register (37,6) Value: %h\n", GRF37_6_buffer[clk]);
        end
        if (GRF37_7_buffer[clk] != GRF37_7_buffer[!clk]) begin
          $fwrite(f, "Register (37,7) Value: %h\n", GRF37_7_buffer[clk]);
        end
        if (GRF37_8_buffer[clk] != GRF37_8_buffer[!clk]) begin
          $fwrite(f, "Register (37,8) Value: %h\n", GRF37_8_buffer[clk]);
        end
        if (GRF37_9_buffer[clk] != GRF37_9_buffer[!clk]) begin
          $fwrite(f, "Register (37,9) Value: %h\n", GRF37_9_buffer[clk]);
        end
        if (GRF37_10_buffer[clk] != GRF37_10_buffer[!clk]) begin
          $fwrite(f, "Register (37,10) Value: %h\n", GRF37_10_buffer[clk]);
        end
        if (GRF37_11_buffer[clk] != GRF37_11_buffer[!clk]) begin
          $fwrite(f, "Register (37,11) Value: %h\n", GRF37_11_buffer[clk]);
        end
        if (GRF37_12_buffer[clk] != GRF37_12_buffer[!clk]) begin
          $fwrite(f, "Register (37,12) Value: %h\n", GRF37_12_buffer[clk]);
        end
        if (GRF37_13_buffer[clk] != GRF37_13_buffer[!clk]) begin
          $fwrite(f, "Register (37,13) Value: %h\n", GRF37_13_buffer[clk]);
        end
        if (GRF37_14_buffer[clk] != GRF37_14_buffer[!clk]) begin
          $fwrite(f, "Register (37,14) Value: %h\n", GRF37_14_buffer[clk]);
        end
        if (GRF37_15_buffer[clk] != GRF37_15_buffer[!clk]) begin
          $fwrite(f, "Register (37,15) Value: %h\n", GRF37_15_buffer[clk]);
        end
        if (GRF37_16_buffer[clk] != GRF37_16_buffer[!clk]) begin
          $fwrite(f, "Register (37,16) Value: %h\n", GRF37_16_buffer[clk]);
        end
        if (GRF37_17_buffer[clk] != GRF37_17_buffer[!clk]) begin
          $fwrite(f, "Register (37,17) Value: %h\n", GRF37_17_buffer[clk]);
        end
        if (GRF37_18_buffer[clk] != GRF37_18_buffer[!clk]) begin
          $fwrite(f, "Register (37,18) Value: %h\n", GRF37_18_buffer[clk]);
        end
        if (GRF37_19_buffer[clk] != GRF37_19_buffer[!clk]) begin
          $fwrite(f, "Register (37,19) Value: %h\n", GRF37_19_buffer[clk]);
        end
        if (GRF37_20_buffer[clk] != GRF37_20_buffer[!clk]) begin
          $fwrite(f, "Register (37,20) Value: %h\n", GRF37_20_buffer[clk]);
        end
        if (GRF37_21_buffer[clk] != GRF37_21_buffer[!clk]) begin
          $fwrite(f, "Register (37,21) Value: %h\n", GRF37_21_buffer[clk]);
        end
        if (GRF37_22_buffer[clk] != GRF37_22_buffer[!clk]) begin
          $fwrite(f, "Register (37,22) Value: %h\n", GRF37_22_buffer[clk]);
        end
        if (GRF37_23_buffer[clk] != GRF37_23_buffer[!clk]) begin
          $fwrite(f, "Register (37,23) Value: %h\n", GRF37_23_buffer[clk]);
        end
        if (GRF37_24_buffer[clk] != GRF37_24_buffer[!clk]) begin
          $fwrite(f, "Register (37,24) Value: %h\n", GRF37_24_buffer[clk]);
        end
        if (GRF37_25_buffer[clk] != GRF37_25_buffer[!clk]) begin
          $fwrite(f, "Register (37,25) Value: %h\n", GRF37_25_buffer[clk]);
        end
        if (GRF37_26_buffer[clk] != GRF37_26_buffer[!clk]) begin
          $fwrite(f, "Register (37,26) Value: %h\n", GRF37_26_buffer[clk]);
        end
        if (GRF37_27_buffer[clk] != GRF37_27_buffer[!clk]) begin
          $fwrite(f, "Register (37,27) Value: %h\n", GRF37_27_buffer[clk]);
        end
        if (GRF37_28_buffer[clk] != GRF37_28_buffer[!clk]) begin
          $fwrite(f, "Register (37,28) Value: %h\n", GRF37_28_buffer[clk]);
        end
        if (GRF37_29_buffer[clk] != GRF37_29_buffer[!clk]) begin
          $fwrite(f, "Register (37,29) Value: %h\n", GRF37_29_buffer[clk]);
        end
        if (GRF37_30_buffer[clk] != GRF37_30_buffer[!clk]) begin
          $fwrite(f, "Register (37,30) Value: %h\n", GRF37_30_buffer[clk]);
        end
        if (GRF37_31_buffer[clk] != GRF37_31_buffer[!clk]) begin
          $fwrite(f, "Register (37,31) Value: %h\n", GRF37_31_buffer[clk]);
        end
        if (GRF38_0_buffer[clk] != GRF38_0_buffer[!clk]) begin
          $fwrite(f, "Register (38,0) Value: %h\n", GRF38_0_buffer[clk]);
        end
        if (GRF38_1_buffer[clk] != GRF38_1_buffer[!clk]) begin
          $fwrite(f, "Register (38,1) Value: %h\n", GRF38_1_buffer[clk]);
        end
        if (GRF38_2_buffer[clk] != GRF38_2_buffer[!clk]) begin
          $fwrite(f, "Register (38,2) Value: %h\n", GRF38_2_buffer[clk]);
        end
        if (GRF38_3_buffer[clk] != GRF38_3_buffer[!clk]) begin
          $fwrite(f, "Register (38,3) Value: %h\n", GRF38_3_buffer[clk]);
        end
        if (GRF38_4_buffer[clk] != GRF38_4_buffer[!clk]) begin
          $fwrite(f, "Register (38,4) Value: %h\n", GRF38_4_buffer[clk]);
        end
        if (GRF38_5_buffer[clk] != GRF38_5_buffer[!clk]) begin
          $fwrite(f, "Register (38,5) Value: %h\n", GRF38_5_buffer[clk]);
        end
        if (GRF38_6_buffer[clk] != GRF38_6_buffer[!clk]) begin
          $fwrite(f, "Register (38,6) Value: %h\n", GRF38_6_buffer[clk]);
        end
        if (GRF38_7_buffer[clk] != GRF38_7_buffer[!clk]) begin
          $fwrite(f, "Register (38,7) Value: %h\n", GRF38_7_buffer[clk]);
        end
        if (GRF38_8_buffer[clk] != GRF38_8_buffer[!clk]) begin
          $fwrite(f, "Register (38,8) Value: %h\n", GRF38_8_buffer[clk]);
        end
        if (GRF38_9_buffer[clk] != GRF38_9_buffer[!clk]) begin
          $fwrite(f, "Register (38,9) Value: %h\n", GRF38_9_buffer[clk]);
        end
        if (GRF38_10_buffer[clk] != GRF38_10_buffer[!clk]) begin
          $fwrite(f, "Register (38,10) Value: %h\n", GRF38_10_buffer[clk]);
        end
        if (GRF38_11_buffer[clk] != GRF38_11_buffer[!clk]) begin
          $fwrite(f, "Register (38,11) Value: %h\n", GRF38_11_buffer[clk]);
        end
        if (GRF38_12_buffer[clk] != GRF38_12_buffer[!clk]) begin
          $fwrite(f, "Register (38,12) Value: %h\n", GRF38_12_buffer[clk]);
        end
        if (GRF38_13_buffer[clk] != GRF38_13_buffer[!clk]) begin
          $fwrite(f, "Register (38,13) Value: %h\n", GRF38_13_buffer[clk]);
        end
        if (GRF38_14_buffer[clk] != GRF38_14_buffer[!clk]) begin
          $fwrite(f, "Register (38,14) Value: %h\n", GRF38_14_buffer[clk]);
        end
        if (GRF38_15_buffer[clk] != GRF38_15_buffer[!clk]) begin
          $fwrite(f, "Register (38,15) Value: %h\n", GRF38_15_buffer[clk]);
        end
        if (GRF38_16_buffer[clk] != GRF38_16_buffer[!clk]) begin
          $fwrite(f, "Register (38,16) Value: %h\n", GRF38_16_buffer[clk]);
        end
        if (GRF38_17_buffer[clk] != GRF38_17_buffer[!clk]) begin
          $fwrite(f, "Register (38,17) Value: %h\n", GRF38_17_buffer[clk]);
        end
        if (GRF38_18_buffer[clk] != GRF38_18_buffer[!clk]) begin
          $fwrite(f, "Register (38,18) Value: %h\n", GRF38_18_buffer[clk]);
        end
        if (GRF38_19_buffer[clk] != GRF38_19_buffer[!clk]) begin
          $fwrite(f, "Register (38,19) Value: %h\n", GRF38_19_buffer[clk]);
        end
        if (GRF38_20_buffer[clk] != GRF38_20_buffer[!clk]) begin
          $fwrite(f, "Register (38,20) Value: %h\n", GRF38_20_buffer[clk]);
        end
        if (GRF38_21_buffer[clk] != GRF38_21_buffer[!clk]) begin
          $fwrite(f, "Register (38,21) Value: %h\n", GRF38_21_buffer[clk]);
        end
        if (GRF38_22_buffer[clk] != GRF38_22_buffer[!clk]) begin
          $fwrite(f, "Register (38,22) Value: %h\n", GRF38_22_buffer[clk]);
        end
        if (GRF38_23_buffer[clk] != GRF38_23_buffer[!clk]) begin
          $fwrite(f, "Register (38,23) Value: %h\n", GRF38_23_buffer[clk]);
        end
        if (GRF38_24_buffer[clk] != GRF38_24_buffer[!clk]) begin
          $fwrite(f, "Register (38,24) Value: %h\n", GRF38_24_buffer[clk]);
        end
        if (GRF38_25_buffer[clk] != GRF38_25_buffer[!clk]) begin
          $fwrite(f, "Register (38,25) Value: %h\n", GRF38_25_buffer[clk]);
        end
        if (GRF38_26_buffer[clk] != GRF38_26_buffer[!clk]) begin
          $fwrite(f, "Register (38,26) Value: %h\n", GRF38_26_buffer[clk]);
        end
        if (GRF38_27_buffer[clk] != GRF38_27_buffer[!clk]) begin
          $fwrite(f, "Register (38,27) Value: %h\n", GRF38_27_buffer[clk]);
        end
        if (GRF38_28_buffer[clk] != GRF38_28_buffer[!clk]) begin
          $fwrite(f, "Register (38,28) Value: %h\n", GRF38_28_buffer[clk]);
        end
        if (GRF38_29_buffer[clk] != GRF38_29_buffer[!clk]) begin
          $fwrite(f, "Register (38,29) Value: %h\n", GRF38_29_buffer[clk]);
        end
        if (GRF38_30_buffer[clk] != GRF38_30_buffer[!clk]) begin
          $fwrite(f, "Register (38,30) Value: %h\n", GRF38_30_buffer[clk]);
        end
        if (GRF38_31_buffer[clk] != GRF38_31_buffer[!clk]) begin
          $fwrite(f, "Register (38,31) Value: %h\n", GRF38_31_buffer[clk]);
        end
        if (GRF39_0_buffer[clk] != GRF39_0_buffer[!clk]) begin
          $fwrite(f, "Register (39,0) Value: %h\n", GRF39_0_buffer[clk]);
        end
        if (GRF39_1_buffer[clk] != GRF39_1_buffer[!clk]) begin
          $fwrite(f, "Register (39,1) Value: %h\n", GRF39_1_buffer[clk]);
        end
        if (GRF39_2_buffer[clk] != GRF39_2_buffer[!clk]) begin
          $fwrite(f, "Register (39,2) Value: %h\n", GRF39_2_buffer[clk]);
        end
        if (GRF39_3_buffer[clk] != GRF39_3_buffer[!clk]) begin
          $fwrite(f, "Register (39,3) Value: %h\n", GRF39_3_buffer[clk]);
        end
        if (GRF39_4_buffer[clk] != GRF39_4_buffer[!clk]) begin
          $fwrite(f, "Register (39,4) Value: %h\n", GRF39_4_buffer[clk]);
        end
        if (GRF39_5_buffer[clk] != GRF39_5_buffer[!clk]) begin
          $fwrite(f, "Register (39,5) Value: %h\n", GRF39_5_buffer[clk]);
        end
        if (GRF39_6_buffer[clk] != GRF39_6_buffer[!clk]) begin
          $fwrite(f, "Register (39,6) Value: %h\n", GRF39_6_buffer[clk]);
        end
        if (GRF39_7_buffer[clk] != GRF39_7_buffer[!clk]) begin
          $fwrite(f, "Register (39,7) Value: %h\n", GRF39_7_buffer[clk]);
        end
        if (GRF39_8_buffer[clk] != GRF39_8_buffer[!clk]) begin
          $fwrite(f, "Register (39,8) Value: %h\n", GRF39_8_buffer[clk]);
        end
        if (GRF39_9_buffer[clk] != GRF39_9_buffer[!clk]) begin
          $fwrite(f, "Register (39,9) Value: %h\n", GRF39_9_buffer[clk]);
        end
        if (GRF39_10_buffer[clk] != GRF39_10_buffer[!clk]) begin
          $fwrite(f, "Register (39,10) Value: %h\n", GRF39_10_buffer[clk]);
        end
        if (GRF39_11_buffer[clk] != GRF39_11_buffer[!clk]) begin
          $fwrite(f, "Register (39,11) Value: %h\n", GRF39_11_buffer[clk]);
        end
        if (GRF39_12_buffer[clk] != GRF39_12_buffer[!clk]) begin
          $fwrite(f, "Register (39,12) Value: %h\n", GRF39_12_buffer[clk]);
        end
        if (GRF39_13_buffer[clk] != GRF39_13_buffer[!clk]) begin
          $fwrite(f, "Register (39,13) Value: %h\n", GRF39_13_buffer[clk]);
        end
        if (GRF39_14_buffer[clk] != GRF39_14_buffer[!clk]) begin
          $fwrite(f, "Register (39,14) Value: %h\n", GRF39_14_buffer[clk]);
        end
        if (GRF39_15_buffer[clk] != GRF39_15_buffer[!clk]) begin
          $fwrite(f, "Register (39,15) Value: %h\n", GRF39_15_buffer[clk]);
        end
        if (GRF39_16_buffer[clk] != GRF39_16_buffer[!clk]) begin
          $fwrite(f, "Register (39,16) Value: %h\n", GRF39_16_buffer[clk]);
        end
        if (GRF39_17_buffer[clk] != GRF39_17_buffer[!clk]) begin
          $fwrite(f, "Register (39,17) Value: %h\n", GRF39_17_buffer[clk]);
        end
        if (GRF39_18_buffer[clk] != GRF39_18_buffer[!clk]) begin
          $fwrite(f, "Register (39,18) Value: %h\n", GRF39_18_buffer[clk]);
        end
        if (GRF39_19_buffer[clk] != GRF39_19_buffer[!clk]) begin
          $fwrite(f, "Register (39,19) Value: %h\n", GRF39_19_buffer[clk]);
        end
        if (GRF39_20_buffer[clk] != GRF39_20_buffer[!clk]) begin
          $fwrite(f, "Register (39,20) Value: %h\n", GRF39_20_buffer[clk]);
        end
        if (GRF39_21_buffer[clk] != GRF39_21_buffer[!clk]) begin
          $fwrite(f, "Register (39,21) Value: %h\n", GRF39_21_buffer[clk]);
        end
        if (GRF39_22_buffer[clk] != GRF39_22_buffer[!clk]) begin
          $fwrite(f, "Register (39,22) Value: %h\n", GRF39_22_buffer[clk]);
        end
        if (GRF39_23_buffer[clk] != GRF39_23_buffer[!clk]) begin
          $fwrite(f, "Register (39,23) Value: %h\n", GRF39_23_buffer[clk]);
        end
        if (GRF39_24_buffer[clk] != GRF39_24_buffer[!clk]) begin
          $fwrite(f, "Register (39,24) Value: %h\n", GRF39_24_buffer[clk]);
        end
        if (GRF39_25_buffer[clk] != GRF39_25_buffer[!clk]) begin
          $fwrite(f, "Register (39,25) Value: %h\n", GRF39_25_buffer[clk]);
        end
        if (GRF39_26_buffer[clk] != GRF39_26_buffer[!clk]) begin
          $fwrite(f, "Register (39,26) Value: %h\n", GRF39_26_buffer[clk]);
        end
        if (GRF39_27_buffer[clk] != GRF39_27_buffer[!clk]) begin
          $fwrite(f, "Register (39,27) Value: %h\n", GRF39_27_buffer[clk]);
        end
        if (GRF39_28_buffer[clk] != GRF39_28_buffer[!clk]) begin
          $fwrite(f, "Register (39,28) Value: %h\n", GRF39_28_buffer[clk]);
        end
        if (GRF39_29_buffer[clk] != GRF39_29_buffer[!clk]) begin
          $fwrite(f, "Register (39,29) Value: %h\n", GRF39_29_buffer[clk]);
        end
        if (GRF39_30_buffer[clk] != GRF39_30_buffer[!clk]) begin
          $fwrite(f, "Register (39,30) Value: %h\n", GRF39_30_buffer[clk]);
        end
        if (GRF39_31_buffer[clk] != GRF39_31_buffer[!clk]) begin
          $fwrite(f, "Register (39,31) Value: %h\n", GRF39_31_buffer[clk]);
        end
        if (GRF40_0_buffer[clk] != GRF40_0_buffer[!clk]) begin
          $fwrite(f, "Register (40,0) Value: %h\n", GRF40_0_buffer[clk]);
        end
        if (GRF40_1_buffer[clk] != GRF40_1_buffer[!clk]) begin
          $fwrite(f, "Register (40,1) Value: %h\n", GRF40_1_buffer[clk]);
        end
        if (GRF40_2_buffer[clk] != GRF40_2_buffer[!clk]) begin
          $fwrite(f, "Register (40,2) Value: %h\n", GRF40_2_buffer[clk]);
        end
        if (GRF40_3_buffer[clk] != GRF40_3_buffer[!clk]) begin
          $fwrite(f, "Register (40,3) Value: %h\n", GRF40_3_buffer[clk]);
        end
        if (GRF40_4_buffer[clk] != GRF40_4_buffer[!clk]) begin
          $fwrite(f, "Register (40,4) Value: %h\n", GRF40_4_buffer[clk]);
        end
        if (GRF40_5_buffer[clk] != GRF40_5_buffer[!clk]) begin
          $fwrite(f, "Register (40,5) Value: %h\n", GRF40_5_buffer[clk]);
        end
        if (GRF40_6_buffer[clk] != GRF40_6_buffer[!clk]) begin
          $fwrite(f, "Register (40,6) Value: %h\n", GRF40_6_buffer[clk]);
        end
        if (GRF40_7_buffer[clk] != GRF40_7_buffer[!clk]) begin
          $fwrite(f, "Register (40,7) Value: %h\n", GRF40_7_buffer[clk]);
        end
        if (GRF40_8_buffer[clk] != GRF40_8_buffer[!clk]) begin
          $fwrite(f, "Register (40,8) Value: %h\n", GRF40_8_buffer[clk]);
        end
        if (GRF40_9_buffer[clk] != GRF40_9_buffer[!clk]) begin
          $fwrite(f, "Register (40,9) Value: %h\n", GRF40_9_buffer[clk]);
        end
        if (GRF40_10_buffer[clk] != GRF40_10_buffer[!clk]) begin
          $fwrite(f, "Register (40,10) Value: %h\n", GRF40_10_buffer[clk]);
        end
        if (GRF40_11_buffer[clk] != GRF40_11_buffer[!clk]) begin
          $fwrite(f, "Register (40,11) Value: %h\n", GRF40_11_buffer[clk]);
        end
        if (GRF40_12_buffer[clk] != GRF40_12_buffer[!clk]) begin
          $fwrite(f, "Register (40,12) Value: %h\n", GRF40_12_buffer[clk]);
        end
        if (GRF40_13_buffer[clk] != GRF40_13_buffer[!clk]) begin
          $fwrite(f, "Register (40,13) Value: %h\n", GRF40_13_buffer[clk]);
        end
        if (GRF40_14_buffer[clk] != GRF40_14_buffer[!clk]) begin
          $fwrite(f, "Register (40,14) Value: %h\n", GRF40_14_buffer[clk]);
        end
        if (GRF40_15_buffer[clk] != GRF40_15_buffer[!clk]) begin
          $fwrite(f, "Register (40,15) Value: %h\n", GRF40_15_buffer[clk]);
        end
        if (GRF40_16_buffer[clk] != GRF40_16_buffer[!clk]) begin
          $fwrite(f, "Register (40,16) Value: %h\n", GRF40_16_buffer[clk]);
        end
        if (GRF40_17_buffer[clk] != GRF40_17_buffer[!clk]) begin
          $fwrite(f, "Register (40,17) Value: %h\n", GRF40_17_buffer[clk]);
        end
        if (GRF40_18_buffer[clk] != GRF40_18_buffer[!clk]) begin
          $fwrite(f, "Register (40,18) Value: %h\n", GRF40_18_buffer[clk]);
        end
        if (GRF40_19_buffer[clk] != GRF40_19_buffer[!clk]) begin
          $fwrite(f, "Register (40,19) Value: %h\n", GRF40_19_buffer[clk]);
        end
        if (GRF40_20_buffer[clk] != GRF40_20_buffer[!clk]) begin
          $fwrite(f, "Register (40,20) Value: %h\n", GRF40_20_buffer[clk]);
        end
        if (GRF40_21_buffer[clk] != GRF40_21_buffer[!clk]) begin
          $fwrite(f, "Register (40,21) Value: %h\n", GRF40_21_buffer[clk]);
        end
        if (GRF40_22_buffer[clk] != GRF40_22_buffer[!clk]) begin
          $fwrite(f, "Register (40,22) Value: %h\n", GRF40_22_buffer[clk]);
        end
        if (GRF40_23_buffer[clk] != GRF40_23_buffer[!clk]) begin
          $fwrite(f, "Register (40,23) Value: %h\n", GRF40_23_buffer[clk]);
        end
        if (GRF40_24_buffer[clk] != GRF40_24_buffer[!clk]) begin
          $fwrite(f, "Register (40,24) Value: %h\n", GRF40_24_buffer[clk]);
        end
        if (GRF40_25_buffer[clk] != GRF40_25_buffer[!clk]) begin
          $fwrite(f, "Register (40,25) Value: %h\n", GRF40_25_buffer[clk]);
        end
        if (GRF40_26_buffer[clk] != GRF40_26_buffer[!clk]) begin
          $fwrite(f, "Register (40,26) Value: %h\n", GRF40_26_buffer[clk]);
        end
        if (GRF40_27_buffer[clk] != GRF40_27_buffer[!clk]) begin
          $fwrite(f, "Register (40,27) Value: %h\n", GRF40_27_buffer[clk]);
        end
        if (GRF40_28_buffer[clk] != GRF40_28_buffer[!clk]) begin
          $fwrite(f, "Register (40,28) Value: %h\n", GRF40_28_buffer[clk]);
        end
        if (GRF40_29_buffer[clk] != GRF40_29_buffer[!clk]) begin
          $fwrite(f, "Register (40,29) Value: %h\n", GRF40_29_buffer[clk]);
        end
        if (GRF40_30_buffer[clk] != GRF40_30_buffer[!clk]) begin
          $fwrite(f, "Register (40,30) Value: %h\n", GRF40_30_buffer[clk]);
        end
        if (GRF40_31_buffer[clk] != GRF40_31_buffer[!clk]) begin
          $fwrite(f, "Register (40,31) Value: %h\n", GRF40_31_buffer[clk]);
        end
        if (GRF41_0_buffer[clk] != GRF41_0_buffer[!clk]) begin
          $fwrite(f, "Register (41,0) Value: %h\n", GRF41_0_buffer[clk]);
        end
        if (GRF41_1_buffer[clk] != GRF41_1_buffer[!clk]) begin
          $fwrite(f, "Register (41,1) Value: %h\n", GRF41_1_buffer[clk]);
        end
        if (GRF41_2_buffer[clk] != GRF41_2_buffer[!clk]) begin
          $fwrite(f, "Register (41,2) Value: %h\n", GRF41_2_buffer[clk]);
        end
        if (GRF41_3_buffer[clk] != GRF41_3_buffer[!clk]) begin
          $fwrite(f, "Register (41,3) Value: %h\n", GRF41_3_buffer[clk]);
        end
        if (GRF41_4_buffer[clk] != GRF41_4_buffer[!clk]) begin
          $fwrite(f, "Register (41,4) Value: %h\n", GRF41_4_buffer[clk]);
        end
        if (GRF41_5_buffer[clk] != GRF41_5_buffer[!clk]) begin
          $fwrite(f, "Register (41,5) Value: %h\n", GRF41_5_buffer[clk]);
        end
        if (GRF41_6_buffer[clk] != GRF41_6_buffer[!clk]) begin
          $fwrite(f, "Register (41,6) Value: %h\n", GRF41_6_buffer[clk]);
        end
        if (GRF41_7_buffer[clk] != GRF41_7_buffer[!clk]) begin
          $fwrite(f, "Register (41,7) Value: %h\n", GRF41_7_buffer[clk]);
        end
        if (GRF41_8_buffer[clk] != GRF41_8_buffer[!clk]) begin
          $fwrite(f, "Register (41,8) Value: %h\n", GRF41_8_buffer[clk]);
        end
        if (GRF41_9_buffer[clk] != GRF41_9_buffer[!clk]) begin
          $fwrite(f, "Register (41,9) Value: %h\n", GRF41_9_buffer[clk]);
        end
        if (GRF41_10_buffer[clk] != GRF41_10_buffer[!clk]) begin
          $fwrite(f, "Register (41,10) Value: %h\n", GRF41_10_buffer[clk]);
        end
        if (GRF41_11_buffer[clk] != GRF41_11_buffer[!clk]) begin
          $fwrite(f, "Register (41,11) Value: %h\n", GRF41_11_buffer[clk]);
        end
        if (GRF41_12_buffer[clk] != GRF41_12_buffer[!clk]) begin
          $fwrite(f, "Register (41,12) Value: %h\n", GRF41_12_buffer[clk]);
        end
        if (GRF41_13_buffer[clk] != GRF41_13_buffer[!clk]) begin
          $fwrite(f, "Register (41,13) Value: %h\n", GRF41_13_buffer[clk]);
        end
        if (GRF41_14_buffer[clk] != GRF41_14_buffer[!clk]) begin
          $fwrite(f, "Register (41,14) Value: %h\n", GRF41_14_buffer[clk]);
        end
        if (GRF41_15_buffer[clk] != GRF41_15_buffer[!clk]) begin
          $fwrite(f, "Register (41,15) Value: %h\n", GRF41_15_buffer[clk]);
        end
        if (GRF41_16_buffer[clk] != GRF41_16_buffer[!clk]) begin
          $fwrite(f, "Register (41,16) Value: %h\n", GRF41_16_buffer[clk]);
        end
        if (GRF41_17_buffer[clk] != GRF41_17_buffer[!clk]) begin
          $fwrite(f, "Register (41,17) Value: %h\n", GRF41_17_buffer[clk]);
        end
        if (GRF41_18_buffer[clk] != GRF41_18_buffer[!clk]) begin
          $fwrite(f, "Register (41,18) Value: %h\n", GRF41_18_buffer[clk]);
        end
        if (GRF41_19_buffer[clk] != GRF41_19_buffer[!clk]) begin
          $fwrite(f, "Register (41,19) Value: %h\n", GRF41_19_buffer[clk]);
        end
        if (GRF41_20_buffer[clk] != GRF41_20_buffer[!clk]) begin
          $fwrite(f, "Register (41,20) Value: %h\n", GRF41_20_buffer[clk]);
        end
        if (GRF41_21_buffer[clk] != GRF41_21_buffer[!clk]) begin
          $fwrite(f, "Register (41,21) Value: %h\n", GRF41_21_buffer[clk]);
        end
        if (GRF41_22_buffer[clk] != GRF41_22_buffer[!clk]) begin
          $fwrite(f, "Register (41,22) Value: %h\n", GRF41_22_buffer[clk]);
        end
        if (GRF41_23_buffer[clk] != GRF41_23_buffer[!clk]) begin
          $fwrite(f, "Register (41,23) Value: %h\n", GRF41_23_buffer[clk]);
        end
        if (GRF41_24_buffer[clk] != GRF41_24_buffer[!clk]) begin
          $fwrite(f, "Register (41,24) Value: %h\n", GRF41_24_buffer[clk]);
        end
        if (GRF41_25_buffer[clk] != GRF41_25_buffer[!clk]) begin
          $fwrite(f, "Register (41,25) Value: %h\n", GRF41_25_buffer[clk]);
        end
        if (GRF41_26_buffer[clk] != GRF41_26_buffer[!clk]) begin
          $fwrite(f, "Register (41,26) Value: %h\n", GRF41_26_buffer[clk]);
        end
        if (GRF41_27_buffer[clk] != GRF41_27_buffer[!clk]) begin
          $fwrite(f, "Register (41,27) Value: %h\n", GRF41_27_buffer[clk]);
        end
        if (GRF41_28_buffer[clk] != GRF41_28_buffer[!clk]) begin
          $fwrite(f, "Register (41,28) Value: %h\n", GRF41_28_buffer[clk]);
        end
        if (GRF41_29_buffer[clk] != GRF41_29_buffer[!clk]) begin
          $fwrite(f, "Register (41,29) Value: %h\n", GRF41_29_buffer[clk]);
        end
        if (GRF41_30_buffer[clk] != GRF41_30_buffer[!clk]) begin
          $fwrite(f, "Register (41,30) Value: %h\n", GRF41_30_buffer[clk]);
        end
        if (GRF41_31_buffer[clk] != GRF41_31_buffer[!clk]) begin
          $fwrite(f, "Register (41,31) Value: %h\n", GRF41_31_buffer[clk]);
        end
        if (GRF42_0_buffer[clk] != GRF42_0_buffer[!clk]) begin
          $fwrite(f, "Register (42,0) Value: %h\n", GRF42_0_buffer[clk]);
        end
        if (GRF42_1_buffer[clk] != GRF42_1_buffer[!clk]) begin
          $fwrite(f, "Register (42,1) Value: %h\n", GRF42_1_buffer[clk]);
        end
        if (GRF42_2_buffer[clk] != GRF42_2_buffer[!clk]) begin
          $fwrite(f, "Register (42,2) Value: %h\n", GRF42_2_buffer[clk]);
        end
        if (GRF42_3_buffer[clk] != GRF42_3_buffer[!clk]) begin
          $fwrite(f, "Register (42,3) Value: %h\n", GRF42_3_buffer[clk]);
        end
        if (GRF42_4_buffer[clk] != GRF42_4_buffer[!clk]) begin
          $fwrite(f, "Register (42,4) Value: %h\n", GRF42_4_buffer[clk]);
        end
        if (GRF42_5_buffer[clk] != GRF42_5_buffer[!clk]) begin
          $fwrite(f, "Register (42,5) Value: %h\n", GRF42_5_buffer[clk]);
        end
        if (GRF42_6_buffer[clk] != GRF42_6_buffer[!clk]) begin
          $fwrite(f, "Register (42,6) Value: %h\n", GRF42_6_buffer[clk]);
        end
        if (GRF42_7_buffer[clk] != GRF42_7_buffer[!clk]) begin
          $fwrite(f, "Register (42,7) Value: %h\n", GRF42_7_buffer[clk]);
        end
        if (GRF42_8_buffer[clk] != GRF42_8_buffer[!clk]) begin
          $fwrite(f, "Register (42,8) Value: %h\n", GRF42_8_buffer[clk]);
        end
        if (GRF42_9_buffer[clk] != GRF42_9_buffer[!clk]) begin
          $fwrite(f, "Register (42,9) Value: %h\n", GRF42_9_buffer[clk]);
        end
        if (GRF42_10_buffer[clk] != GRF42_10_buffer[!clk]) begin
          $fwrite(f, "Register (42,10) Value: %h\n", GRF42_10_buffer[clk]);
        end
        if (GRF42_11_buffer[clk] != GRF42_11_buffer[!clk]) begin
          $fwrite(f, "Register (42,11) Value: %h\n", GRF42_11_buffer[clk]);
        end
        if (GRF42_12_buffer[clk] != GRF42_12_buffer[!clk]) begin
          $fwrite(f, "Register (42,12) Value: %h\n", GRF42_12_buffer[clk]);
        end
        if (GRF42_13_buffer[clk] != GRF42_13_buffer[!clk]) begin
          $fwrite(f, "Register (42,13) Value: %h\n", GRF42_13_buffer[clk]);
        end
        if (GRF42_14_buffer[clk] != GRF42_14_buffer[!clk]) begin
          $fwrite(f, "Register (42,14) Value: %h\n", GRF42_14_buffer[clk]);
        end
        if (GRF42_15_buffer[clk] != GRF42_15_buffer[!clk]) begin
          $fwrite(f, "Register (42,15) Value: %h\n", GRF42_15_buffer[clk]);
        end
        if (GRF42_16_buffer[clk] != GRF42_16_buffer[!clk]) begin
          $fwrite(f, "Register (42,16) Value: %h\n", GRF42_16_buffer[clk]);
        end
        if (GRF42_17_buffer[clk] != GRF42_17_buffer[!clk]) begin
          $fwrite(f, "Register (42,17) Value: %h\n", GRF42_17_buffer[clk]);
        end
        if (GRF42_18_buffer[clk] != GRF42_18_buffer[!clk]) begin
          $fwrite(f, "Register (42,18) Value: %h\n", GRF42_18_buffer[clk]);
        end
        if (GRF42_19_buffer[clk] != GRF42_19_buffer[!clk]) begin
          $fwrite(f, "Register (42,19) Value: %h\n", GRF42_19_buffer[clk]);
        end
        if (GRF42_20_buffer[clk] != GRF42_20_buffer[!clk]) begin
          $fwrite(f, "Register (42,20) Value: %h\n", GRF42_20_buffer[clk]);
        end
        if (GRF42_21_buffer[clk] != GRF42_21_buffer[!clk]) begin
          $fwrite(f, "Register (42,21) Value: %h\n", GRF42_21_buffer[clk]);
        end
        if (GRF42_22_buffer[clk] != GRF42_22_buffer[!clk]) begin
          $fwrite(f, "Register (42,22) Value: %h\n", GRF42_22_buffer[clk]);
        end
        if (GRF42_23_buffer[clk] != GRF42_23_buffer[!clk]) begin
          $fwrite(f, "Register (42,23) Value: %h\n", GRF42_23_buffer[clk]);
        end
        if (GRF42_24_buffer[clk] != GRF42_24_buffer[!clk]) begin
          $fwrite(f, "Register (42,24) Value: %h\n", GRF42_24_buffer[clk]);
        end
        if (GRF42_25_buffer[clk] != GRF42_25_buffer[!clk]) begin
          $fwrite(f, "Register (42,25) Value: %h\n", GRF42_25_buffer[clk]);
        end
        if (GRF42_26_buffer[clk] != GRF42_26_buffer[!clk]) begin
          $fwrite(f, "Register (42,26) Value: %h\n", GRF42_26_buffer[clk]);
        end
        if (GRF42_27_buffer[clk] != GRF42_27_buffer[!clk]) begin
          $fwrite(f, "Register (42,27) Value: %h\n", GRF42_27_buffer[clk]);
        end
        if (GRF42_28_buffer[clk] != GRF42_28_buffer[!clk]) begin
          $fwrite(f, "Register (42,28) Value: %h\n", GRF42_28_buffer[clk]);
        end
        if (GRF42_29_buffer[clk] != GRF42_29_buffer[!clk]) begin
          $fwrite(f, "Register (42,29) Value: %h\n", GRF42_29_buffer[clk]);
        end
        if (GRF42_30_buffer[clk] != GRF42_30_buffer[!clk]) begin
          $fwrite(f, "Register (42,30) Value: %h\n", GRF42_30_buffer[clk]);
        end
        if (GRF42_31_buffer[clk] != GRF42_31_buffer[!clk]) begin
          $fwrite(f, "Register (42,31) Value: %h\n", GRF42_31_buffer[clk]);
        end
        if (GRF43_0_buffer[clk] != GRF43_0_buffer[!clk]) begin
          $fwrite(f, "Register (43,0) Value: %h\n", GRF43_0_buffer[clk]);
        end
        if (GRF43_1_buffer[clk] != GRF43_1_buffer[!clk]) begin
          $fwrite(f, "Register (43,1) Value: %h\n", GRF43_1_buffer[clk]);
        end
        if (GRF43_2_buffer[clk] != GRF43_2_buffer[!clk]) begin
          $fwrite(f, "Register (43,2) Value: %h\n", GRF43_2_buffer[clk]);
        end
        if (GRF43_3_buffer[clk] != GRF43_3_buffer[!clk]) begin
          $fwrite(f, "Register (43,3) Value: %h\n", GRF43_3_buffer[clk]);
        end
        if (GRF43_4_buffer[clk] != GRF43_4_buffer[!clk]) begin
          $fwrite(f, "Register (43,4) Value: %h\n", GRF43_4_buffer[clk]);
        end
        if (GRF43_5_buffer[clk] != GRF43_5_buffer[!clk]) begin
          $fwrite(f, "Register (43,5) Value: %h\n", GRF43_5_buffer[clk]);
        end
        if (GRF43_6_buffer[clk] != GRF43_6_buffer[!clk]) begin
          $fwrite(f, "Register (43,6) Value: %h\n", GRF43_6_buffer[clk]);
        end
        if (GRF43_7_buffer[clk] != GRF43_7_buffer[!clk]) begin
          $fwrite(f, "Register (43,7) Value: %h\n", GRF43_7_buffer[clk]);
        end
        if (GRF43_8_buffer[clk] != GRF43_8_buffer[!clk]) begin
          $fwrite(f, "Register (43,8) Value: %h\n", GRF43_8_buffer[clk]);
        end
        if (GRF43_9_buffer[clk] != GRF43_9_buffer[!clk]) begin
          $fwrite(f, "Register (43,9) Value: %h\n", GRF43_9_buffer[clk]);
        end
        if (GRF43_10_buffer[clk] != GRF43_10_buffer[!clk]) begin
          $fwrite(f, "Register (43,10) Value: %h\n", GRF43_10_buffer[clk]);
        end
        if (GRF43_11_buffer[clk] != GRF43_11_buffer[!clk]) begin
          $fwrite(f, "Register (43,11) Value: %h\n", GRF43_11_buffer[clk]);
        end
        if (GRF43_12_buffer[clk] != GRF43_12_buffer[!clk]) begin
          $fwrite(f, "Register (43,12) Value: %h\n", GRF43_12_buffer[clk]);
        end
        if (GRF43_13_buffer[clk] != GRF43_13_buffer[!clk]) begin
          $fwrite(f, "Register (43,13) Value: %h\n", GRF43_13_buffer[clk]);
        end
        if (GRF43_14_buffer[clk] != GRF43_14_buffer[!clk]) begin
          $fwrite(f, "Register (43,14) Value: %h\n", GRF43_14_buffer[clk]);
        end
        if (GRF43_15_buffer[clk] != GRF43_15_buffer[!clk]) begin
          $fwrite(f, "Register (43,15) Value: %h\n", GRF43_15_buffer[clk]);
        end
        if (GRF43_16_buffer[clk] != GRF43_16_buffer[!clk]) begin
          $fwrite(f, "Register (43,16) Value: %h\n", GRF43_16_buffer[clk]);
        end
        if (GRF43_17_buffer[clk] != GRF43_17_buffer[!clk]) begin
          $fwrite(f, "Register (43,17) Value: %h\n", GRF43_17_buffer[clk]);
        end
        if (GRF43_18_buffer[clk] != GRF43_18_buffer[!clk]) begin
          $fwrite(f, "Register (43,18) Value: %h\n", GRF43_18_buffer[clk]);
        end
        if (GRF43_19_buffer[clk] != GRF43_19_buffer[!clk]) begin
          $fwrite(f, "Register (43,19) Value: %h\n", GRF43_19_buffer[clk]);
        end
        if (GRF43_20_buffer[clk] != GRF43_20_buffer[!clk]) begin
          $fwrite(f, "Register (43,20) Value: %h\n", GRF43_20_buffer[clk]);
        end
        if (GRF43_21_buffer[clk] != GRF43_21_buffer[!clk]) begin
          $fwrite(f, "Register (43,21) Value: %h\n", GRF43_21_buffer[clk]);
        end
        if (GRF43_22_buffer[clk] != GRF43_22_buffer[!clk]) begin
          $fwrite(f, "Register (43,22) Value: %h\n", GRF43_22_buffer[clk]);
        end
        if (GRF43_23_buffer[clk] != GRF43_23_buffer[!clk]) begin
          $fwrite(f, "Register (43,23) Value: %h\n", GRF43_23_buffer[clk]);
        end
        if (GRF43_24_buffer[clk] != GRF43_24_buffer[!clk]) begin
          $fwrite(f, "Register (43,24) Value: %h\n", GRF43_24_buffer[clk]);
        end
        if (GRF43_25_buffer[clk] != GRF43_25_buffer[!clk]) begin
          $fwrite(f, "Register (43,25) Value: %h\n", GRF43_25_buffer[clk]);
        end
        if (GRF43_26_buffer[clk] != GRF43_26_buffer[!clk]) begin
          $fwrite(f, "Register (43,26) Value: %h\n", GRF43_26_buffer[clk]);
        end
        if (GRF43_27_buffer[clk] != GRF43_27_buffer[!clk]) begin
          $fwrite(f, "Register (43,27) Value: %h\n", GRF43_27_buffer[clk]);
        end
        if (GRF43_28_buffer[clk] != GRF43_28_buffer[!clk]) begin
          $fwrite(f, "Register (43,28) Value: %h\n", GRF43_28_buffer[clk]);
        end
        if (GRF43_29_buffer[clk] != GRF43_29_buffer[!clk]) begin
          $fwrite(f, "Register (43,29) Value: %h\n", GRF43_29_buffer[clk]);
        end
        if (GRF43_30_buffer[clk] != GRF43_30_buffer[!clk]) begin
          $fwrite(f, "Register (43,30) Value: %h\n", GRF43_30_buffer[clk]);
        end
        if (GRF43_31_buffer[clk] != GRF43_31_buffer[!clk]) begin
          $fwrite(f, "Register (43,31) Value: %h\n", GRF43_31_buffer[clk]);
        end
        if (GRF44_0_buffer[clk] != GRF44_0_buffer[!clk]) begin
          $fwrite(f, "Register (44,0) Value: %h\n", GRF44_0_buffer[clk]);
        end
        if (GRF44_1_buffer[clk] != GRF44_1_buffer[!clk]) begin
          $fwrite(f, "Register (44,1) Value: %h\n", GRF44_1_buffer[clk]);
        end
        if (GRF44_2_buffer[clk] != GRF44_2_buffer[!clk]) begin
          $fwrite(f, "Register (44,2) Value: %h\n", GRF44_2_buffer[clk]);
        end
        if (GRF44_3_buffer[clk] != GRF44_3_buffer[!clk]) begin
          $fwrite(f, "Register (44,3) Value: %h\n", GRF44_3_buffer[clk]);
        end
        if (GRF44_4_buffer[clk] != GRF44_4_buffer[!clk]) begin
          $fwrite(f, "Register (44,4) Value: %h\n", GRF44_4_buffer[clk]);
        end
        if (GRF44_5_buffer[clk] != GRF44_5_buffer[!clk]) begin
          $fwrite(f, "Register (44,5) Value: %h\n", GRF44_5_buffer[clk]);
        end
        if (GRF44_6_buffer[clk] != GRF44_6_buffer[!clk]) begin
          $fwrite(f, "Register (44,6) Value: %h\n", GRF44_6_buffer[clk]);
        end
        if (GRF44_7_buffer[clk] != GRF44_7_buffer[!clk]) begin
          $fwrite(f, "Register (44,7) Value: %h\n", GRF44_7_buffer[clk]);
        end
        if (GRF44_8_buffer[clk] != GRF44_8_buffer[!clk]) begin
          $fwrite(f, "Register (44,8) Value: %h\n", GRF44_8_buffer[clk]);
        end
        if (GRF44_9_buffer[clk] != GRF44_9_buffer[!clk]) begin
          $fwrite(f, "Register (44,9) Value: %h\n", GRF44_9_buffer[clk]);
        end
        if (GRF44_10_buffer[clk] != GRF44_10_buffer[!clk]) begin
          $fwrite(f, "Register (44,10) Value: %h\n", GRF44_10_buffer[clk]);
        end
        if (GRF44_11_buffer[clk] != GRF44_11_buffer[!clk]) begin
          $fwrite(f, "Register (44,11) Value: %h\n", GRF44_11_buffer[clk]);
        end
        if (GRF44_12_buffer[clk] != GRF44_12_buffer[!clk]) begin
          $fwrite(f, "Register (44,12) Value: %h\n", GRF44_12_buffer[clk]);
        end
        if (GRF44_13_buffer[clk] != GRF44_13_buffer[!clk]) begin
          $fwrite(f, "Register (44,13) Value: %h\n", GRF44_13_buffer[clk]);
        end
        if (GRF44_14_buffer[clk] != GRF44_14_buffer[!clk]) begin
          $fwrite(f, "Register (44,14) Value: %h\n", GRF44_14_buffer[clk]);
        end
        if (GRF44_15_buffer[clk] != GRF44_15_buffer[!clk]) begin
          $fwrite(f, "Register (44,15) Value: %h\n", GRF44_15_buffer[clk]);
        end
        if (GRF44_16_buffer[clk] != GRF44_16_buffer[!clk]) begin
          $fwrite(f, "Register (44,16) Value: %h\n", GRF44_16_buffer[clk]);
        end
        if (GRF44_17_buffer[clk] != GRF44_17_buffer[!clk]) begin
          $fwrite(f, "Register (44,17) Value: %h\n", GRF44_17_buffer[clk]);
        end
        if (GRF44_18_buffer[clk] != GRF44_18_buffer[!clk]) begin
          $fwrite(f, "Register (44,18) Value: %h\n", GRF44_18_buffer[clk]);
        end
        if (GRF44_19_buffer[clk] != GRF44_19_buffer[!clk]) begin
          $fwrite(f, "Register (44,19) Value: %h\n", GRF44_19_buffer[clk]);
        end
        if (GRF44_20_buffer[clk] != GRF44_20_buffer[!clk]) begin
          $fwrite(f, "Register (44,20) Value: %h\n", GRF44_20_buffer[clk]);
        end
        if (GRF44_21_buffer[clk] != GRF44_21_buffer[!clk]) begin
          $fwrite(f, "Register (44,21) Value: %h\n", GRF44_21_buffer[clk]);
        end
        if (GRF44_22_buffer[clk] != GRF44_22_buffer[!clk]) begin
          $fwrite(f, "Register (44,22) Value: %h\n", GRF44_22_buffer[clk]);
        end
        if (GRF44_23_buffer[clk] != GRF44_23_buffer[!clk]) begin
          $fwrite(f, "Register (44,23) Value: %h\n", GRF44_23_buffer[clk]);
        end
        if (GRF44_24_buffer[clk] != GRF44_24_buffer[!clk]) begin
          $fwrite(f, "Register (44,24) Value: %h\n", GRF44_24_buffer[clk]);
        end
        if (GRF44_25_buffer[clk] != GRF44_25_buffer[!clk]) begin
          $fwrite(f, "Register (44,25) Value: %h\n", GRF44_25_buffer[clk]);
        end
        if (GRF44_26_buffer[clk] != GRF44_26_buffer[!clk]) begin
          $fwrite(f, "Register (44,26) Value: %h\n", GRF44_26_buffer[clk]);
        end
        if (GRF44_27_buffer[clk] != GRF44_27_buffer[!clk]) begin
          $fwrite(f, "Register (44,27) Value: %h\n", GRF44_27_buffer[clk]);
        end
        if (GRF44_28_buffer[clk] != GRF44_28_buffer[!clk]) begin
          $fwrite(f, "Register (44,28) Value: %h\n", GRF44_28_buffer[clk]);
        end
        if (GRF44_29_buffer[clk] != GRF44_29_buffer[!clk]) begin
          $fwrite(f, "Register (44,29) Value: %h\n", GRF44_29_buffer[clk]);
        end
        if (GRF44_30_buffer[clk] != GRF44_30_buffer[!clk]) begin
          $fwrite(f, "Register (44,30) Value: %h\n", GRF44_30_buffer[clk]);
        end
        if (GRF44_31_buffer[clk] != GRF44_31_buffer[!clk]) begin
          $fwrite(f, "Register (44,31) Value: %h\n", GRF44_31_buffer[clk]);
        end
        if (GRF45_0_buffer[clk] != GRF45_0_buffer[!clk]) begin
          $fwrite(f, "Register (45,0) Value: %h\n", GRF45_0_buffer[clk]);
        end
        if (GRF45_1_buffer[clk] != GRF45_1_buffer[!clk]) begin
          $fwrite(f, "Register (45,1) Value: %h\n", GRF45_1_buffer[clk]);
        end
        if (GRF45_2_buffer[clk] != GRF45_2_buffer[!clk]) begin
          $fwrite(f, "Register (45,2) Value: %h\n", GRF45_2_buffer[clk]);
        end
        if (GRF45_3_buffer[clk] != GRF45_3_buffer[!clk]) begin
          $fwrite(f, "Register (45,3) Value: %h\n", GRF45_3_buffer[clk]);
        end
        if (GRF45_4_buffer[clk] != GRF45_4_buffer[!clk]) begin
          $fwrite(f, "Register (45,4) Value: %h\n", GRF45_4_buffer[clk]);
        end
        if (GRF45_5_buffer[clk] != GRF45_5_buffer[!clk]) begin
          $fwrite(f, "Register (45,5) Value: %h\n", GRF45_5_buffer[clk]);
        end
        if (GRF45_6_buffer[clk] != GRF45_6_buffer[!clk]) begin
          $fwrite(f, "Register (45,6) Value: %h\n", GRF45_6_buffer[clk]);
        end
        if (GRF45_7_buffer[clk] != GRF45_7_buffer[!clk]) begin
          $fwrite(f, "Register (45,7) Value: %h\n", GRF45_7_buffer[clk]);
        end
        if (GRF45_8_buffer[clk] != GRF45_8_buffer[!clk]) begin
          $fwrite(f, "Register (45,8) Value: %h\n", GRF45_8_buffer[clk]);
        end
        if (GRF45_9_buffer[clk] != GRF45_9_buffer[!clk]) begin
          $fwrite(f, "Register (45,9) Value: %h\n", GRF45_9_buffer[clk]);
        end
        if (GRF45_10_buffer[clk] != GRF45_10_buffer[!clk]) begin
          $fwrite(f, "Register (45,10) Value: %h\n", GRF45_10_buffer[clk]);
        end
        if (GRF45_11_buffer[clk] != GRF45_11_buffer[!clk]) begin
          $fwrite(f, "Register (45,11) Value: %h\n", GRF45_11_buffer[clk]);
        end
        if (GRF45_12_buffer[clk] != GRF45_12_buffer[!clk]) begin
          $fwrite(f, "Register (45,12) Value: %h\n", GRF45_12_buffer[clk]);
        end
        if (GRF45_13_buffer[clk] != GRF45_13_buffer[!clk]) begin
          $fwrite(f, "Register (45,13) Value: %h\n", GRF45_13_buffer[clk]);
        end
        if (GRF45_14_buffer[clk] != GRF45_14_buffer[!clk]) begin
          $fwrite(f, "Register (45,14) Value: %h\n", GRF45_14_buffer[clk]);
        end
        if (GRF45_15_buffer[clk] != GRF45_15_buffer[!clk]) begin
          $fwrite(f, "Register (45,15) Value: %h\n", GRF45_15_buffer[clk]);
        end
        if (GRF45_16_buffer[clk] != GRF45_16_buffer[!clk]) begin
          $fwrite(f, "Register (45,16) Value: %h\n", GRF45_16_buffer[clk]);
        end
        if (GRF45_17_buffer[clk] != GRF45_17_buffer[!clk]) begin
          $fwrite(f, "Register (45,17) Value: %h\n", GRF45_17_buffer[clk]);
        end
        if (GRF45_18_buffer[clk] != GRF45_18_buffer[!clk]) begin
          $fwrite(f, "Register (45,18) Value: %h\n", GRF45_18_buffer[clk]);
        end
        if (GRF45_19_buffer[clk] != GRF45_19_buffer[!clk]) begin
          $fwrite(f, "Register (45,19) Value: %h\n", GRF45_19_buffer[clk]);
        end
        if (GRF45_20_buffer[clk] != GRF45_20_buffer[!clk]) begin
          $fwrite(f, "Register (45,20) Value: %h\n", GRF45_20_buffer[clk]);
        end
        if (GRF45_21_buffer[clk] != GRF45_21_buffer[!clk]) begin
          $fwrite(f, "Register (45,21) Value: %h\n", GRF45_21_buffer[clk]);
        end
        if (GRF45_22_buffer[clk] != GRF45_22_buffer[!clk]) begin
          $fwrite(f, "Register (45,22) Value: %h\n", GRF45_22_buffer[clk]);
        end
        if (GRF45_23_buffer[clk] != GRF45_23_buffer[!clk]) begin
          $fwrite(f, "Register (45,23) Value: %h\n", GRF45_23_buffer[clk]);
        end
        if (GRF45_24_buffer[clk] != GRF45_24_buffer[!clk]) begin
          $fwrite(f, "Register (45,24) Value: %h\n", GRF45_24_buffer[clk]);
        end
        if (GRF45_25_buffer[clk] != GRF45_25_buffer[!clk]) begin
          $fwrite(f, "Register (45,25) Value: %h\n", GRF45_25_buffer[clk]);
        end
        if (GRF45_26_buffer[clk] != GRF45_26_buffer[!clk]) begin
          $fwrite(f, "Register (45,26) Value: %h\n", GRF45_26_buffer[clk]);
        end
        if (GRF45_27_buffer[clk] != GRF45_27_buffer[!clk]) begin
          $fwrite(f, "Register (45,27) Value: %h\n", GRF45_27_buffer[clk]);
        end
        if (GRF45_28_buffer[clk] != GRF45_28_buffer[!clk]) begin
          $fwrite(f, "Register (45,28) Value: %h\n", GRF45_28_buffer[clk]);
        end
        if (GRF45_29_buffer[clk] != GRF45_29_buffer[!clk]) begin
          $fwrite(f, "Register (45,29) Value: %h\n", GRF45_29_buffer[clk]);
        end
        if (GRF45_30_buffer[clk] != GRF45_30_buffer[!clk]) begin
          $fwrite(f, "Register (45,30) Value: %h\n", GRF45_30_buffer[clk]);
        end
        if (GRF45_31_buffer[clk] != GRF45_31_buffer[!clk]) begin
          $fwrite(f, "Register (45,31) Value: %h\n", GRF45_31_buffer[clk]);
        end
        if (GRF46_0_buffer[clk] != GRF46_0_buffer[!clk]) begin
          $fwrite(f, "Register (46,0) Value: %h\n", GRF46_0_buffer[clk]);
        end
        if (GRF46_1_buffer[clk] != GRF46_1_buffer[!clk]) begin
          $fwrite(f, "Register (46,1) Value: %h\n", GRF46_1_buffer[clk]);
        end
        if (GRF46_2_buffer[clk] != GRF46_2_buffer[!clk]) begin
          $fwrite(f, "Register (46,2) Value: %h\n", GRF46_2_buffer[clk]);
        end
        if (GRF46_3_buffer[clk] != GRF46_3_buffer[!clk]) begin
          $fwrite(f, "Register (46,3) Value: %h\n", GRF46_3_buffer[clk]);
        end
        if (GRF46_4_buffer[clk] != GRF46_4_buffer[!clk]) begin
          $fwrite(f, "Register (46,4) Value: %h\n", GRF46_4_buffer[clk]);
        end
        if (GRF46_5_buffer[clk] != GRF46_5_buffer[!clk]) begin
          $fwrite(f, "Register (46,5) Value: %h\n", GRF46_5_buffer[clk]);
        end
        if (GRF46_6_buffer[clk] != GRF46_6_buffer[!clk]) begin
          $fwrite(f, "Register (46,6) Value: %h\n", GRF46_6_buffer[clk]);
        end
        if (GRF46_7_buffer[clk] != GRF46_7_buffer[!clk]) begin
          $fwrite(f, "Register (46,7) Value: %h\n", GRF46_7_buffer[clk]);
        end
        if (GRF46_8_buffer[clk] != GRF46_8_buffer[!clk]) begin
          $fwrite(f, "Register (46,8) Value: %h\n", GRF46_8_buffer[clk]);
        end
        if (GRF46_9_buffer[clk] != GRF46_9_buffer[!clk]) begin
          $fwrite(f, "Register (46,9) Value: %h\n", GRF46_9_buffer[clk]);
        end
        if (GRF46_10_buffer[clk] != GRF46_10_buffer[!clk]) begin
          $fwrite(f, "Register (46,10) Value: %h\n", GRF46_10_buffer[clk]);
        end
        if (GRF46_11_buffer[clk] != GRF46_11_buffer[!clk]) begin
          $fwrite(f, "Register (46,11) Value: %h\n", GRF46_11_buffer[clk]);
        end
        if (GRF46_12_buffer[clk] != GRF46_12_buffer[!clk]) begin
          $fwrite(f, "Register (46,12) Value: %h\n", GRF46_12_buffer[clk]);
        end
        if (GRF46_13_buffer[clk] != GRF46_13_buffer[!clk]) begin
          $fwrite(f, "Register (46,13) Value: %h\n", GRF46_13_buffer[clk]);
        end
        if (GRF46_14_buffer[clk] != GRF46_14_buffer[!clk]) begin
          $fwrite(f, "Register (46,14) Value: %h\n", GRF46_14_buffer[clk]);
        end
        if (GRF46_15_buffer[clk] != GRF46_15_buffer[!clk]) begin
          $fwrite(f, "Register (46,15) Value: %h\n", GRF46_15_buffer[clk]);
        end
        if (GRF46_16_buffer[clk] != GRF46_16_buffer[!clk]) begin
          $fwrite(f, "Register (46,16) Value: %h\n", GRF46_16_buffer[clk]);
        end
        if (GRF46_17_buffer[clk] != GRF46_17_buffer[!clk]) begin
          $fwrite(f, "Register (46,17) Value: %h\n", GRF46_17_buffer[clk]);
        end
        if (GRF46_18_buffer[clk] != GRF46_18_buffer[!clk]) begin
          $fwrite(f, "Register (46,18) Value: %h\n", GRF46_18_buffer[clk]);
        end
        if (GRF46_19_buffer[clk] != GRF46_19_buffer[!clk]) begin
          $fwrite(f, "Register (46,19) Value: %h\n", GRF46_19_buffer[clk]);
        end
        if (GRF46_20_buffer[clk] != GRF46_20_buffer[!clk]) begin
          $fwrite(f, "Register (46,20) Value: %h\n", GRF46_20_buffer[clk]);
        end
        if (GRF46_21_buffer[clk] != GRF46_21_buffer[!clk]) begin
          $fwrite(f, "Register (46,21) Value: %h\n", GRF46_21_buffer[clk]);
        end
        if (GRF46_22_buffer[clk] != GRF46_22_buffer[!clk]) begin
          $fwrite(f, "Register (46,22) Value: %h\n", GRF46_22_buffer[clk]);
        end
        if (GRF46_23_buffer[clk] != GRF46_23_buffer[!clk]) begin
          $fwrite(f, "Register (46,23) Value: %h\n", GRF46_23_buffer[clk]);
        end
        if (GRF46_24_buffer[clk] != GRF46_24_buffer[!clk]) begin
          $fwrite(f, "Register (46,24) Value: %h\n", GRF46_24_buffer[clk]);
        end
        if (GRF46_25_buffer[clk] != GRF46_25_buffer[!clk]) begin
          $fwrite(f, "Register (46,25) Value: %h\n", GRF46_25_buffer[clk]);
        end
        if (GRF46_26_buffer[clk] != GRF46_26_buffer[!clk]) begin
          $fwrite(f, "Register (46,26) Value: %h\n", GRF46_26_buffer[clk]);
        end
        if (GRF46_27_buffer[clk] != GRF46_27_buffer[!clk]) begin
          $fwrite(f, "Register (46,27) Value: %h\n", GRF46_27_buffer[clk]);
        end
        if (GRF46_28_buffer[clk] != GRF46_28_buffer[!clk]) begin
          $fwrite(f, "Register (46,28) Value: %h\n", GRF46_28_buffer[clk]);
        end
        if (GRF46_29_buffer[clk] != GRF46_29_buffer[!clk]) begin
          $fwrite(f, "Register (46,29) Value: %h\n", GRF46_29_buffer[clk]);
        end
        if (GRF46_30_buffer[clk] != GRF46_30_buffer[!clk]) begin
          $fwrite(f, "Register (46,30) Value: %h\n", GRF46_30_buffer[clk]);
        end
        if (GRF46_31_buffer[clk] != GRF46_31_buffer[!clk]) begin
          $fwrite(f, "Register (46,31) Value: %h\n", GRF46_31_buffer[clk]);
        end
        if (GRF47_0_buffer[clk] != GRF47_0_buffer[!clk]) begin
          $fwrite(f, "Register (47,0) Value: %h\n", GRF47_0_buffer[clk]);
        end
        if (GRF47_1_buffer[clk] != GRF47_1_buffer[!clk]) begin
          $fwrite(f, "Register (47,1) Value: %h\n", GRF47_1_buffer[clk]);
        end
        if (GRF47_2_buffer[clk] != GRF47_2_buffer[!clk]) begin
          $fwrite(f, "Register (47,2) Value: %h\n", GRF47_2_buffer[clk]);
        end
        if (GRF47_3_buffer[clk] != GRF47_3_buffer[!clk]) begin
          $fwrite(f, "Register (47,3) Value: %h\n", GRF47_3_buffer[clk]);
        end
        if (GRF47_4_buffer[clk] != GRF47_4_buffer[!clk]) begin
          $fwrite(f, "Register (47,4) Value: %h\n", GRF47_4_buffer[clk]);
        end
        if (GRF47_5_buffer[clk] != GRF47_5_buffer[!clk]) begin
          $fwrite(f, "Register (47,5) Value: %h\n", GRF47_5_buffer[clk]);
        end
        if (GRF47_6_buffer[clk] != GRF47_6_buffer[!clk]) begin
          $fwrite(f, "Register (47,6) Value: %h\n", GRF47_6_buffer[clk]);
        end
        if (GRF47_7_buffer[clk] != GRF47_7_buffer[!clk]) begin
          $fwrite(f, "Register (47,7) Value: %h\n", GRF47_7_buffer[clk]);
        end
        if (GRF47_8_buffer[clk] != GRF47_8_buffer[!clk]) begin
          $fwrite(f, "Register (47,8) Value: %h\n", GRF47_8_buffer[clk]);
        end
        if (GRF47_9_buffer[clk] != GRF47_9_buffer[!clk]) begin
          $fwrite(f, "Register (47,9) Value: %h\n", GRF47_9_buffer[clk]);
        end
        if (GRF47_10_buffer[clk] != GRF47_10_buffer[!clk]) begin
          $fwrite(f, "Register (47,10) Value: %h\n", GRF47_10_buffer[clk]);
        end
        if (GRF47_11_buffer[clk] != GRF47_11_buffer[!clk]) begin
          $fwrite(f, "Register (47,11) Value: %h\n", GRF47_11_buffer[clk]);
        end
        if (GRF47_12_buffer[clk] != GRF47_12_buffer[!clk]) begin
          $fwrite(f, "Register (47,12) Value: %h\n", GRF47_12_buffer[clk]);
        end
        if (GRF47_13_buffer[clk] != GRF47_13_buffer[!clk]) begin
          $fwrite(f, "Register (47,13) Value: %h\n", GRF47_13_buffer[clk]);
        end
        if (GRF47_14_buffer[clk] != GRF47_14_buffer[!clk]) begin
          $fwrite(f, "Register (47,14) Value: %h\n", GRF47_14_buffer[clk]);
        end
        if (GRF47_15_buffer[clk] != GRF47_15_buffer[!clk]) begin
          $fwrite(f, "Register (47,15) Value: %h\n", GRF47_15_buffer[clk]);
        end
        if (GRF47_16_buffer[clk] != GRF47_16_buffer[!clk]) begin
          $fwrite(f, "Register (47,16) Value: %h\n", GRF47_16_buffer[clk]);
        end
        if (GRF47_17_buffer[clk] != GRF47_17_buffer[!clk]) begin
          $fwrite(f, "Register (47,17) Value: %h\n", GRF47_17_buffer[clk]);
        end
        if (GRF47_18_buffer[clk] != GRF47_18_buffer[!clk]) begin
          $fwrite(f, "Register (47,18) Value: %h\n", GRF47_18_buffer[clk]);
        end
        if (GRF47_19_buffer[clk] != GRF47_19_buffer[!clk]) begin
          $fwrite(f, "Register (47,19) Value: %h\n", GRF47_19_buffer[clk]);
        end
        if (GRF47_20_buffer[clk] != GRF47_20_buffer[!clk]) begin
          $fwrite(f, "Register (47,20) Value: %h\n", GRF47_20_buffer[clk]);
        end
        if (GRF47_21_buffer[clk] != GRF47_21_buffer[!clk]) begin
          $fwrite(f, "Register (47,21) Value: %h\n", GRF47_21_buffer[clk]);
        end
        if (GRF47_22_buffer[clk] != GRF47_22_buffer[!clk]) begin
          $fwrite(f, "Register (47,22) Value: %h\n", GRF47_22_buffer[clk]);
        end
        if (GRF47_23_buffer[clk] != GRF47_23_buffer[!clk]) begin
          $fwrite(f, "Register (47,23) Value: %h\n", GRF47_23_buffer[clk]);
        end
        if (GRF47_24_buffer[clk] != GRF47_24_buffer[!clk]) begin
          $fwrite(f, "Register (47,24) Value: %h\n", GRF47_24_buffer[clk]);
        end
        if (GRF47_25_buffer[clk] != GRF47_25_buffer[!clk]) begin
          $fwrite(f, "Register (47,25) Value: %h\n", GRF47_25_buffer[clk]);
        end
        if (GRF47_26_buffer[clk] != GRF47_26_buffer[!clk]) begin
          $fwrite(f, "Register (47,26) Value: %h\n", GRF47_26_buffer[clk]);
        end
        if (GRF47_27_buffer[clk] != GRF47_27_buffer[!clk]) begin
          $fwrite(f, "Register (47,27) Value: %h\n", GRF47_27_buffer[clk]);
        end
        if (GRF47_28_buffer[clk] != GRF47_28_buffer[!clk]) begin
          $fwrite(f, "Register (47,28) Value: %h\n", GRF47_28_buffer[clk]);
        end
        if (GRF47_29_buffer[clk] != GRF47_29_buffer[!clk]) begin
          $fwrite(f, "Register (47,29) Value: %h\n", GRF47_29_buffer[clk]);
        end
        if (GRF47_30_buffer[clk] != GRF47_30_buffer[!clk]) begin
          $fwrite(f, "Register (47,30) Value: %h\n", GRF47_30_buffer[clk]);
        end
        if (GRF47_31_buffer[clk] != GRF47_31_buffer[!clk]) begin
          $fwrite(f, "Register (47,31) Value: %h\n", GRF47_31_buffer[clk]);
        end
        if (GRF48_0_buffer[clk] != GRF48_0_buffer[!clk]) begin
          $fwrite(f, "Register (48,0) Value: %h\n", GRF48_0_buffer[clk]);
        end
        if (GRF48_1_buffer[clk] != GRF48_1_buffer[!clk]) begin
          $fwrite(f, "Register (48,1) Value: %h\n", GRF48_1_buffer[clk]);
        end
        if (GRF48_2_buffer[clk] != GRF48_2_buffer[!clk]) begin
          $fwrite(f, "Register (48,2) Value: %h\n", GRF48_2_buffer[clk]);
        end
        if (GRF48_3_buffer[clk] != GRF48_3_buffer[!clk]) begin
          $fwrite(f, "Register (48,3) Value: %h\n", GRF48_3_buffer[clk]);
        end
        if (GRF48_4_buffer[clk] != GRF48_4_buffer[!clk]) begin
          $fwrite(f, "Register (48,4) Value: %h\n", GRF48_4_buffer[clk]);
        end
        if (GRF48_5_buffer[clk] != GRF48_5_buffer[!clk]) begin
          $fwrite(f, "Register (48,5) Value: %h\n", GRF48_5_buffer[clk]);
        end
        if (GRF48_6_buffer[clk] != GRF48_6_buffer[!clk]) begin
          $fwrite(f, "Register (48,6) Value: %h\n", GRF48_6_buffer[clk]);
        end
        if (GRF48_7_buffer[clk] != GRF48_7_buffer[!clk]) begin
          $fwrite(f, "Register (48,7) Value: %h\n", GRF48_7_buffer[clk]);
        end
        if (GRF48_8_buffer[clk] != GRF48_8_buffer[!clk]) begin
          $fwrite(f, "Register (48,8) Value: %h\n", GRF48_8_buffer[clk]);
        end
        if (GRF48_9_buffer[clk] != GRF48_9_buffer[!clk]) begin
          $fwrite(f, "Register (48,9) Value: %h\n", GRF48_9_buffer[clk]);
        end
        if (GRF48_10_buffer[clk] != GRF48_10_buffer[!clk]) begin
          $fwrite(f, "Register (48,10) Value: %h\n", GRF48_10_buffer[clk]);
        end
        if (GRF48_11_buffer[clk] != GRF48_11_buffer[!clk]) begin
          $fwrite(f, "Register (48,11) Value: %h\n", GRF48_11_buffer[clk]);
        end
        if (GRF48_12_buffer[clk] != GRF48_12_buffer[!clk]) begin
          $fwrite(f, "Register (48,12) Value: %h\n", GRF48_12_buffer[clk]);
        end
        if (GRF48_13_buffer[clk] != GRF48_13_buffer[!clk]) begin
          $fwrite(f, "Register (48,13) Value: %h\n", GRF48_13_buffer[clk]);
        end
        if (GRF48_14_buffer[clk] != GRF48_14_buffer[!clk]) begin
          $fwrite(f, "Register (48,14) Value: %h\n", GRF48_14_buffer[clk]);
        end
        if (GRF48_15_buffer[clk] != GRF48_15_buffer[!clk]) begin
          $fwrite(f, "Register (48,15) Value: %h\n", GRF48_15_buffer[clk]);
        end
        if (GRF48_16_buffer[clk] != GRF48_16_buffer[!clk]) begin
          $fwrite(f, "Register (48,16) Value: %h\n", GRF48_16_buffer[clk]);
        end
        if (GRF48_17_buffer[clk] != GRF48_17_buffer[!clk]) begin
          $fwrite(f, "Register (48,17) Value: %h\n", GRF48_17_buffer[clk]);
        end
        if (GRF48_18_buffer[clk] != GRF48_18_buffer[!clk]) begin
          $fwrite(f, "Register (48,18) Value: %h\n", GRF48_18_buffer[clk]);
        end
        if (GRF48_19_buffer[clk] != GRF48_19_buffer[!clk]) begin
          $fwrite(f, "Register (48,19) Value: %h\n", GRF48_19_buffer[clk]);
        end
        if (GRF48_20_buffer[clk] != GRF48_20_buffer[!clk]) begin
          $fwrite(f, "Register (48,20) Value: %h\n", GRF48_20_buffer[clk]);
        end
        if (GRF48_21_buffer[clk] != GRF48_21_buffer[!clk]) begin
          $fwrite(f, "Register (48,21) Value: %h\n", GRF48_21_buffer[clk]);
        end
        if (GRF48_22_buffer[clk] != GRF48_22_buffer[!clk]) begin
          $fwrite(f, "Register (48,22) Value: %h\n", GRF48_22_buffer[clk]);
        end
        if (GRF48_23_buffer[clk] != GRF48_23_buffer[!clk]) begin
          $fwrite(f, "Register (48,23) Value: %h\n", GRF48_23_buffer[clk]);
        end
        if (GRF48_24_buffer[clk] != GRF48_24_buffer[!clk]) begin
          $fwrite(f, "Register (48,24) Value: %h\n", GRF48_24_buffer[clk]);
        end
        if (GRF48_25_buffer[clk] != GRF48_25_buffer[!clk]) begin
          $fwrite(f, "Register (48,25) Value: %h\n", GRF48_25_buffer[clk]);
        end
        if (GRF48_26_buffer[clk] != GRF48_26_buffer[!clk]) begin
          $fwrite(f, "Register (48,26) Value: %h\n", GRF48_26_buffer[clk]);
        end
        if (GRF48_27_buffer[clk] != GRF48_27_buffer[!clk]) begin
          $fwrite(f, "Register (48,27) Value: %h\n", GRF48_27_buffer[clk]);
        end
        if (GRF48_28_buffer[clk] != GRF48_28_buffer[!clk]) begin
          $fwrite(f, "Register (48,28) Value: %h\n", GRF48_28_buffer[clk]);
        end
        if (GRF48_29_buffer[clk] != GRF48_29_buffer[!clk]) begin
          $fwrite(f, "Register (48,29) Value: %h\n", GRF48_29_buffer[clk]);
        end
        if (GRF48_30_buffer[clk] != GRF48_30_buffer[!clk]) begin
          $fwrite(f, "Register (48,30) Value: %h\n", GRF48_30_buffer[clk]);
        end
        if (GRF48_31_buffer[clk] != GRF48_31_buffer[!clk]) begin
          $fwrite(f, "Register (48,31) Value: %h\n", GRF48_31_buffer[clk]);
        end
        if (GRF49_0_buffer[clk] != GRF49_0_buffer[!clk]) begin
          $fwrite(f, "Register (49,0) Value: %h\n", GRF49_0_buffer[clk]);
        end
        if (GRF49_1_buffer[clk] != GRF49_1_buffer[!clk]) begin
          $fwrite(f, "Register (49,1) Value: %h\n", GRF49_1_buffer[clk]);
        end
        if (GRF49_2_buffer[clk] != GRF49_2_buffer[!clk]) begin
          $fwrite(f, "Register (49,2) Value: %h\n", GRF49_2_buffer[clk]);
        end
        if (GRF49_3_buffer[clk] != GRF49_3_buffer[!clk]) begin
          $fwrite(f, "Register (49,3) Value: %h\n", GRF49_3_buffer[clk]);
        end
        if (GRF49_4_buffer[clk] != GRF49_4_buffer[!clk]) begin
          $fwrite(f, "Register (49,4) Value: %h\n", GRF49_4_buffer[clk]);
        end
        if (GRF49_5_buffer[clk] != GRF49_5_buffer[!clk]) begin
          $fwrite(f, "Register (49,5) Value: %h\n", GRF49_5_buffer[clk]);
        end
        if (GRF49_6_buffer[clk] != GRF49_6_buffer[!clk]) begin
          $fwrite(f, "Register (49,6) Value: %h\n", GRF49_6_buffer[clk]);
        end
        if (GRF49_7_buffer[clk] != GRF49_7_buffer[!clk]) begin
          $fwrite(f, "Register (49,7) Value: %h\n", GRF49_7_buffer[clk]);
        end
        if (GRF49_8_buffer[clk] != GRF49_8_buffer[!clk]) begin
          $fwrite(f, "Register (49,8) Value: %h\n", GRF49_8_buffer[clk]);
        end
        if (GRF49_9_buffer[clk] != GRF49_9_buffer[!clk]) begin
          $fwrite(f, "Register (49,9) Value: %h\n", GRF49_9_buffer[clk]);
        end
        if (GRF49_10_buffer[clk] != GRF49_10_buffer[!clk]) begin
          $fwrite(f, "Register (49,10) Value: %h\n", GRF49_10_buffer[clk]);
        end
        if (GRF49_11_buffer[clk] != GRF49_11_buffer[!clk]) begin
          $fwrite(f, "Register (49,11) Value: %h\n", GRF49_11_buffer[clk]);
        end
        if (GRF49_12_buffer[clk] != GRF49_12_buffer[!clk]) begin
          $fwrite(f, "Register (49,12) Value: %h\n", GRF49_12_buffer[clk]);
        end
        if (GRF49_13_buffer[clk] != GRF49_13_buffer[!clk]) begin
          $fwrite(f, "Register (49,13) Value: %h\n", GRF49_13_buffer[clk]);
        end
        if (GRF49_14_buffer[clk] != GRF49_14_buffer[!clk]) begin
          $fwrite(f, "Register (49,14) Value: %h\n", GRF49_14_buffer[clk]);
        end
        if (GRF49_15_buffer[clk] != GRF49_15_buffer[!clk]) begin
          $fwrite(f, "Register (49,15) Value: %h\n", GRF49_15_buffer[clk]);
        end
        if (GRF49_16_buffer[clk] != GRF49_16_buffer[!clk]) begin
          $fwrite(f, "Register (49,16) Value: %h\n", GRF49_16_buffer[clk]);
        end
        if (GRF49_17_buffer[clk] != GRF49_17_buffer[!clk]) begin
          $fwrite(f, "Register (49,17) Value: %h\n", GRF49_17_buffer[clk]);
        end
        if (GRF49_18_buffer[clk] != GRF49_18_buffer[!clk]) begin
          $fwrite(f, "Register (49,18) Value: %h\n", GRF49_18_buffer[clk]);
        end
        if (GRF49_19_buffer[clk] != GRF49_19_buffer[!clk]) begin
          $fwrite(f, "Register (49,19) Value: %h\n", GRF49_19_buffer[clk]);
        end
        if (GRF49_20_buffer[clk] != GRF49_20_buffer[!clk]) begin
          $fwrite(f, "Register (49,20) Value: %h\n", GRF49_20_buffer[clk]);
        end
        if (GRF49_21_buffer[clk] != GRF49_21_buffer[!clk]) begin
          $fwrite(f, "Register (49,21) Value: %h\n", GRF49_21_buffer[clk]);
        end
        if (GRF49_22_buffer[clk] != GRF49_22_buffer[!clk]) begin
          $fwrite(f, "Register (49,22) Value: %h\n", GRF49_22_buffer[clk]);
        end
        if (GRF49_23_buffer[clk] != GRF49_23_buffer[!clk]) begin
          $fwrite(f, "Register (49,23) Value: %h\n", GRF49_23_buffer[clk]);
        end
        if (GRF49_24_buffer[clk] != GRF49_24_buffer[!clk]) begin
          $fwrite(f, "Register (49,24) Value: %h\n", GRF49_24_buffer[clk]);
        end
        if (GRF49_25_buffer[clk] != GRF49_25_buffer[!clk]) begin
          $fwrite(f, "Register (49,25) Value: %h\n", GRF49_25_buffer[clk]);
        end
        if (GRF49_26_buffer[clk] != GRF49_26_buffer[!clk]) begin
          $fwrite(f, "Register (49,26) Value: %h\n", GRF49_26_buffer[clk]);
        end
        if (GRF49_27_buffer[clk] != GRF49_27_buffer[!clk]) begin
          $fwrite(f, "Register (49,27) Value: %h\n", GRF49_27_buffer[clk]);
        end
        if (GRF49_28_buffer[clk] != GRF49_28_buffer[!clk]) begin
          $fwrite(f, "Register (49,28) Value: %h\n", GRF49_28_buffer[clk]);
        end
        if (GRF49_29_buffer[clk] != GRF49_29_buffer[!clk]) begin
          $fwrite(f, "Register (49,29) Value: %h\n", GRF49_29_buffer[clk]);
        end
        if (GRF49_30_buffer[clk] != GRF49_30_buffer[!clk]) begin
          $fwrite(f, "Register (49,30) Value: %h\n", GRF49_30_buffer[clk]);
        end
        if (GRF49_31_buffer[clk] != GRF49_31_buffer[!clk]) begin
          $fwrite(f, "Register (49,31) Value: %h\n", GRF49_31_buffer[clk]);
        end
        if (GRF50_0_buffer[clk] != GRF50_0_buffer[!clk]) begin
          $fwrite(f, "Register (50,0) Value: %h\n", GRF50_0_buffer[clk]);
        end
        if (GRF50_1_buffer[clk] != GRF50_1_buffer[!clk]) begin
          $fwrite(f, "Register (50,1) Value: %h\n", GRF50_1_buffer[clk]);
        end
        if (GRF50_2_buffer[clk] != GRF50_2_buffer[!clk]) begin
          $fwrite(f, "Register (50,2) Value: %h\n", GRF50_2_buffer[clk]);
        end
        if (GRF50_3_buffer[clk] != GRF50_3_buffer[!clk]) begin
          $fwrite(f, "Register (50,3) Value: %h\n", GRF50_3_buffer[clk]);
        end
        if (GRF50_4_buffer[clk] != GRF50_4_buffer[!clk]) begin
          $fwrite(f, "Register (50,4) Value: %h\n", GRF50_4_buffer[clk]);
        end
        if (GRF50_5_buffer[clk] != GRF50_5_buffer[!clk]) begin
          $fwrite(f, "Register (50,5) Value: %h\n", GRF50_5_buffer[clk]);
        end
        if (GRF50_6_buffer[clk] != GRF50_6_buffer[!clk]) begin
          $fwrite(f, "Register (50,6) Value: %h\n", GRF50_6_buffer[clk]);
        end
        if (GRF50_7_buffer[clk] != GRF50_7_buffer[!clk]) begin
          $fwrite(f, "Register (50,7) Value: %h\n", GRF50_7_buffer[clk]);
        end
        if (GRF50_8_buffer[clk] != GRF50_8_buffer[!clk]) begin
          $fwrite(f, "Register (50,8) Value: %h\n", GRF50_8_buffer[clk]);
        end
        if (GRF50_9_buffer[clk] != GRF50_9_buffer[!clk]) begin
          $fwrite(f, "Register (50,9) Value: %h\n", GRF50_9_buffer[clk]);
        end
        if (GRF50_10_buffer[clk] != GRF50_10_buffer[!clk]) begin
          $fwrite(f, "Register (50,10) Value: %h\n", GRF50_10_buffer[clk]);
        end
        if (GRF50_11_buffer[clk] != GRF50_11_buffer[!clk]) begin
          $fwrite(f, "Register (50,11) Value: %h\n", GRF50_11_buffer[clk]);
        end
        if (GRF50_12_buffer[clk] != GRF50_12_buffer[!clk]) begin
          $fwrite(f, "Register (50,12) Value: %h\n", GRF50_12_buffer[clk]);
        end
        if (GRF50_13_buffer[clk] != GRF50_13_buffer[!clk]) begin
          $fwrite(f, "Register (50,13) Value: %h\n", GRF50_13_buffer[clk]);
        end
        if (GRF50_14_buffer[clk] != GRF50_14_buffer[!clk]) begin
          $fwrite(f, "Register (50,14) Value: %h\n", GRF50_14_buffer[clk]);
        end
        if (GRF50_15_buffer[clk] != GRF50_15_buffer[!clk]) begin
          $fwrite(f, "Register (50,15) Value: %h\n", GRF50_15_buffer[clk]);
        end
        if (GRF50_16_buffer[clk] != GRF50_16_buffer[!clk]) begin
          $fwrite(f, "Register (50,16) Value: %h\n", GRF50_16_buffer[clk]);
        end
        if (GRF50_17_buffer[clk] != GRF50_17_buffer[!clk]) begin
          $fwrite(f, "Register (50,17) Value: %h\n", GRF50_17_buffer[clk]);
        end
        if (GRF50_18_buffer[clk] != GRF50_18_buffer[!clk]) begin
          $fwrite(f, "Register (50,18) Value: %h\n", GRF50_18_buffer[clk]);
        end
        if (GRF50_19_buffer[clk] != GRF50_19_buffer[!clk]) begin
          $fwrite(f, "Register (50,19) Value: %h\n", GRF50_19_buffer[clk]);
        end
        if (GRF50_20_buffer[clk] != GRF50_20_buffer[!clk]) begin
          $fwrite(f, "Register (50,20) Value: %h\n", GRF50_20_buffer[clk]);
        end
        if (GRF50_21_buffer[clk] != GRF50_21_buffer[!clk]) begin
          $fwrite(f, "Register (50,21) Value: %h\n", GRF50_21_buffer[clk]);
        end
        if (GRF50_22_buffer[clk] != GRF50_22_buffer[!clk]) begin
          $fwrite(f, "Register (50,22) Value: %h\n", GRF50_22_buffer[clk]);
        end
        if (GRF50_23_buffer[clk] != GRF50_23_buffer[!clk]) begin
          $fwrite(f, "Register (50,23) Value: %h\n", GRF50_23_buffer[clk]);
        end
        if (GRF50_24_buffer[clk] != GRF50_24_buffer[!clk]) begin
          $fwrite(f, "Register (50,24) Value: %h\n", GRF50_24_buffer[clk]);
        end
        if (GRF50_25_buffer[clk] != GRF50_25_buffer[!clk]) begin
          $fwrite(f, "Register (50,25) Value: %h\n", GRF50_25_buffer[clk]);
        end
        if (GRF50_26_buffer[clk] != GRF50_26_buffer[!clk]) begin
          $fwrite(f, "Register (50,26) Value: %h\n", GRF50_26_buffer[clk]);
        end
        if (GRF50_27_buffer[clk] != GRF50_27_buffer[!clk]) begin
          $fwrite(f, "Register (50,27) Value: %h\n", GRF50_27_buffer[clk]);
        end
        if (GRF50_28_buffer[clk] != GRF50_28_buffer[!clk]) begin
          $fwrite(f, "Register (50,28) Value: %h\n", GRF50_28_buffer[clk]);
        end
        if (GRF50_29_buffer[clk] != GRF50_29_buffer[!clk]) begin
          $fwrite(f, "Register (50,29) Value: %h\n", GRF50_29_buffer[clk]);
        end
        if (GRF50_30_buffer[clk] != GRF50_30_buffer[!clk]) begin
          $fwrite(f, "Register (50,30) Value: %h\n", GRF50_30_buffer[clk]);
        end
        if (GRF50_31_buffer[clk] != GRF50_31_buffer[!clk]) begin
          $fwrite(f, "Register (50,31) Value: %h\n", GRF50_31_buffer[clk]);
        end
        if (GRF51_0_buffer[clk] != GRF51_0_buffer[!clk]) begin
          $fwrite(f, "Register (51,0) Value: %h\n", GRF51_0_buffer[clk]);
        end
        if (GRF51_1_buffer[clk] != GRF51_1_buffer[!clk]) begin
          $fwrite(f, "Register (51,1) Value: %h\n", GRF51_1_buffer[clk]);
        end
        if (GRF51_2_buffer[clk] != GRF51_2_buffer[!clk]) begin
          $fwrite(f, "Register (51,2) Value: %h\n", GRF51_2_buffer[clk]);
        end
        if (GRF51_3_buffer[clk] != GRF51_3_buffer[!clk]) begin
          $fwrite(f, "Register (51,3) Value: %h\n", GRF51_3_buffer[clk]);
        end
        if (GRF51_4_buffer[clk] != GRF51_4_buffer[!clk]) begin
          $fwrite(f, "Register (51,4) Value: %h\n", GRF51_4_buffer[clk]);
        end
        if (GRF51_5_buffer[clk] != GRF51_5_buffer[!clk]) begin
          $fwrite(f, "Register (51,5) Value: %h\n", GRF51_5_buffer[clk]);
        end
        if (GRF51_6_buffer[clk] != GRF51_6_buffer[!clk]) begin
          $fwrite(f, "Register (51,6) Value: %h\n", GRF51_6_buffer[clk]);
        end
        if (GRF51_7_buffer[clk] != GRF51_7_buffer[!clk]) begin
          $fwrite(f, "Register (51,7) Value: %h\n", GRF51_7_buffer[clk]);
        end
        if (GRF51_8_buffer[clk] != GRF51_8_buffer[!clk]) begin
          $fwrite(f, "Register (51,8) Value: %h\n", GRF51_8_buffer[clk]);
        end
        if (GRF51_9_buffer[clk] != GRF51_9_buffer[!clk]) begin
          $fwrite(f, "Register (51,9) Value: %h\n", GRF51_9_buffer[clk]);
        end
        if (GRF51_10_buffer[clk] != GRF51_10_buffer[!clk]) begin
          $fwrite(f, "Register (51,10) Value: %h\n", GRF51_10_buffer[clk]);
        end
        if (GRF51_11_buffer[clk] != GRF51_11_buffer[!clk]) begin
          $fwrite(f, "Register (51,11) Value: %h\n", GRF51_11_buffer[clk]);
        end
        if (GRF51_12_buffer[clk] != GRF51_12_buffer[!clk]) begin
          $fwrite(f, "Register (51,12) Value: %h\n", GRF51_12_buffer[clk]);
        end
        if (GRF51_13_buffer[clk] != GRF51_13_buffer[!clk]) begin
          $fwrite(f, "Register (51,13) Value: %h\n", GRF51_13_buffer[clk]);
        end
        if (GRF51_14_buffer[clk] != GRF51_14_buffer[!clk]) begin
          $fwrite(f, "Register (51,14) Value: %h\n", GRF51_14_buffer[clk]);
        end
        if (GRF51_15_buffer[clk] != GRF51_15_buffer[!clk]) begin
          $fwrite(f, "Register (51,15) Value: %h\n", GRF51_15_buffer[clk]);
        end
        if (GRF51_16_buffer[clk] != GRF51_16_buffer[!clk]) begin
          $fwrite(f, "Register (51,16) Value: %h\n", GRF51_16_buffer[clk]);
        end
        if (GRF51_17_buffer[clk] != GRF51_17_buffer[!clk]) begin
          $fwrite(f, "Register (51,17) Value: %h\n", GRF51_17_buffer[clk]);
        end
        if (GRF51_18_buffer[clk] != GRF51_18_buffer[!clk]) begin
          $fwrite(f, "Register (51,18) Value: %h\n", GRF51_18_buffer[clk]);
        end
        if (GRF51_19_buffer[clk] != GRF51_19_buffer[!clk]) begin
          $fwrite(f, "Register (51,19) Value: %h\n", GRF51_19_buffer[clk]);
        end
        if (GRF51_20_buffer[clk] != GRF51_20_buffer[!clk]) begin
          $fwrite(f, "Register (51,20) Value: %h\n", GRF51_20_buffer[clk]);
        end
        if (GRF51_21_buffer[clk] != GRF51_21_buffer[!clk]) begin
          $fwrite(f, "Register (51,21) Value: %h\n", GRF51_21_buffer[clk]);
        end
        if (GRF51_22_buffer[clk] != GRF51_22_buffer[!clk]) begin
          $fwrite(f, "Register (51,22) Value: %h\n", GRF51_22_buffer[clk]);
        end
        if (GRF51_23_buffer[clk] != GRF51_23_buffer[!clk]) begin
          $fwrite(f, "Register (51,23) Value: %h\n", GRF51_23_buffer[clk]);
        end
        if (GRF51_24_buffer[clk] != GRF51_24_buffer[!clk]) begin
          $fwrite(f, "Register (51,24) Value: %h\n", GRF51_24_buffer[clk]);
        end
        if (GRF51_25_buffer[clk] != GRF51_25_buffer[!clk]) begin
          $fwrite(f, "Register (51,25) Value: %h\n", GRF51_25_buffer[clk]);
        end
        if (GRF51_26_buffer[clk] != GRF51_26_buffer[!clk]) begin
          $fwrite(f, "Register (51,26) Value: %h\n", GRF51_26_buffer[clk]);
        end
        if (GRF51_27_buffer[clk] != GRF51_27_buffer[!clk]) begin
          $fwrite(f, "Register (51,27) Value: %h\n", GRF51_27_buffer[clk]);
        end
        if (GRF51_28_buffer[clk] != GRF51_28_buffer[!clk]) begin
          $fwrite(f, "Register (51,28) Value: %h\n", GRF51_28_buffer[clk]);
        end
        if (GRF51_29_buffer[clk] != GRF51_29_buffer[!clk]) begin
          $fwrite(f, "Register (51,29) Value: %h\n", GRF51_29_buffer[clk]);
        end
        if (GRF51_30_buffer[clk] != GRF51_30_buffer[!clk]) begin
          $fwrite(f, "Register (51,30) Value: %h\n", GRF51_30_buffer[clk]);
        end
        if (GRF51_31_buffer[clk] != GRF51_31_buffer[!clk]) begin
          $fwrite(f, "Register (51,31) Value: %h\n", GRF51_31_buffer[clk]);
        end
        if (GRF52_0_buffer[clk] != GRF52_0_buffer[!clk]) begin
          $fwrite(f, "Register (52,0) Value: %h\n", GRF52_0_buffer[clk]);
        end
        if (GRF52_1_buffer[clk] != GRF52_1_buffer[!clk]) begin
          $fwrite(f, "Register (52,1) Value: %h\n", GRF52_1_buffer[clk]);
        end
        if (GRF52_2_buffer[clk] != GRF52_2_buffer[!clk]) begin
          $fwrite(f, "Register (52,2) Value: %h\n", GRF52_2_buffer[clk]);
        end
        if (GRF52_3_buffer[clk] != GRF52_3_buffer[!clk]) begin
          $fwrite(f, "Register (52,3) Value: %h\n", GRF52_3_buffer[clk]);
        end
        if (GRF52_4_buffer[clk] != GRF52_4_buffer[!clk]) begin
          $fwrite(f, "Register (52,4) Value: %h\n", GRF52_4_buffer[clk]);
        end
        if (GRF52_5_buffer[clk] != GRF52_5_buffer[!clk]) begin
          $fwrite(f, "Register (52,5) Value: %h\n", GRF52_5_buffer[clk]);
        end
        if (GRF52_6_buffer[clk] != GRF52_6_buffer[!clk]) begin
          $fwrite(f, "Register (52,6) Value: %h\n", GRF52_6_buffer[clk]);
        end
        if (GRF52_7_buffer[clk] != GRF52_7_buffer[!clk]) begin
          $fwrite(f, "Register (52,7) Value: %h\n", GRF52_7_buffer[clk]);
        end
        if (GRF52_8_buffer[clk] != GRF52_8_buffer[!clk]) begin
          $fwrite(f, "Register (52,8) Value: %h\n", GRF52_8_buffer[clk]);
        end
        if (GRF52_9_buffer[clk] != GRF52_9_buffer[!clk]) begin
          $fwrite(f, "Register (52,9) Value: %h\n", GRF52_9_buffer[clk]);
        end
        if (GRF52_10_buffer[clk] != GRF52_10_buffer[!clk]) begin
          $fwrite(f, "Register (52,10) Value: %h\n", GRF52_10_buffer[clk]);
        end
        if (GRF52_11_buffer[clk] != GRF52_11_buffer[!clk]) begin
          $fwrite(f, "Register (52,11) Value: %h\n", GRF52_11_buffer[clk]);
        end
        if (GRF52_12_buffer[clk] != GRF52_12_buffer[!clk]) begin
          $fwrite(f, "Register (52,12) Value: %h\n", GRF52_12_buffer[clk]);
        end
        if (GRF52_13_buffer[clk] != GRF52_13_buffer[!clk]) begin
          $fwrite(f, "Register (52,13) Value: %h\n", GRF52_13_buffer[clk]);
        end
        if (GRF52_14_buffer[clk] != GRF52_14_buffer[!clk]) begin
          $fwrite(f, "Register (52,14) Value: %h\n", GRF52_14_buffer[clk]);
        end
        if (GRF52_15_buffer[clk] != GRF52_15_buffer[!clk]) begin
          $fwrite(f, "Register (52,15) Value: %h\n", GRF52_15_buffer[clk]);
        end
        if (GRF52_16_buffer[clk] != GRF52_16_buffer[!clk]) begin
          $fwrite(f, "Register (52,16) Value: %h\n", GRF52_16_buffer[clk]);
        end
        if (GRF52_17_buffer[clk] != GRF52_17_buffer[!clk]) begin
          $fwrite(f, "Register (52,17) Value: %h\n", GRF52_17_buffer[clk]);
        end
        if (GRF52_18_buffer[clk] != GRF52_18_buffer[!clk]) begin
          $fwrite(f, "Register (52,18) Value: %h\n", GRF52_18_buffer[clk]);
        end
        if (GRF52_19_buffer[clk] != GRF52_19_buffer[!clk]) begin
          $fwrite(f, "Register (52,19) Value: %h\n", GRF52_19_buffer[clk]);
        end
        if (GRF52_20_buffer[clk] != GRF52_20_buffer[!clk]) begin
          $fwrite(f, "Register (52,20) Value: %h\n", GRF52_20_buffer[clk]);
        end
        if (GRF52_21_buffer[clk] != GRF52_21_buffer[!clk]) begin
          $fwrite(f, "Register (52,21) Value: %h\n", GRF52_21_buffer[clk]);
        end
        if (GRF52_22_buffer[clk] != GRF52_22_buffer[!clk]) begin
          $fwrite(f, "Register (52,22) Value: %h\n", GRF52_22_buffer[clk]);
        end
        if (GRF52_23_buffer[clk] != GRF52_23_buffer[!clk]) begin
          $fwrite(f, "Register (52,23) Value: %h\n", GRF52_23_buffer[clk]);
        end
        if (GRF52_24_buffer[clk] != GRF52_24_buffer[!clk]) begin
          $fwrite(f, "Register (52,24) Value: %h\n", GRF52_24_buffer[clk]);
        end
        if (GRF52_25_buffer[clk] != GRF52_25_buffer[!clk]) begin
          $fwrite(f, "Register (52,25) Value: %h\n", GRF52_25_buffer[clk]);
        end
        if (GRF52_26_buffer[clk] != GRF52_26_buffer[!clk]) begin
          $fwrite(f, "Register (52,26) Value: %h\n", GRF52_26_buffer[clk]);
        end
        if (GRF52_27_buffer[clk] != GRF52_27_buffer[!clk]) begin
          $fwrite(f, "Register (52,27) Value: %h\n", GRF52_27_buffer[clk]);
        end
        if (GRF52_28_buffer[clk] != GRF52_28_buffer[!clk]) begin
          $fwrite(f, "Register (52,28) Value: %h\n", GRF52_28_buffer[clk]);
        end
        if (GRF52_29_buffer[clk] != GRF52_29_buffer[!clk]) begin
          $fwrite(f, "Register (52,29) Value: %h\n", GRF52_29_buffer[clk]);
        end
        if (GRF52_30_buffer[clk] != GRF52_30_buffer[!clk]) begin
          $fwrite(f, "Register (52,30) Value: %h\n", GRF52_30_buffer[clk]);
        end
        if (GRF52_31_buffer[clk] != GRF52_31_buffer[!clk]) begin
          $fwrite(f, "Register (52,31) Value: %h\n", GRF52_31_buffer[clk]);
        end
        if (GRF53_0_buffer[clk] != GRF53_0_buffer[!clk]) begin
          $fwrite(f, "Register (53,0) Value: %h\n", GRF53_0_buffer[clk]);
        end
        if (GRF53_1_buffer[clk] != GRF53_1_buffer[!clk]) begin
          $fwrite(f, "Register (53,1) Value: %h\n", GRF53_1_buffer[clk]);
        end
        if (GRF53_2_buffer[clk] != GRF53_2_buffer[!clk]) begin
          $fwrite(f, "Register (53,2) Value: %h\n", GRF53_2_buffer[clk]);
        end
        if (GRF53_3_buffer[clk] != GRF53_3_buffer[!clk]) begin
          $fwrite(f, "Register (53,3) Value: %h\n", GRF53_3_buffer[clk]);
        end
        if (GRF53_4_buffer[clk] != GRF53_4_buffer[!clk]) begin
          $fwrite(f, "Register (53,4) Value: %h\n", GRF53_4_buffer[clk]);
        end
        if (GRF53_5_buffer[clk] != GRF53_5_buffer[!clk]) begin
          $fwrite(f, "Register (53,5) Value: %h\n", GRF53_5_buffer[clk]);
        end
        if (GRF53_6_buffer[clk] != GRF53_6_buffer[!clk]) begin
          $fwrite(f, "Register (53,6) Value: %h\n", GRF53_6_buffer[clk]);
        end
        if (GRF53_7_buffer[clk] != GRF53_7_buffer[!clk]) begin
          $fwrite(f, "Register (53,7) Value: %h\n", GRF53_7_buffer[clk]);
        end
        if (GRF53_8_buffer[clk] != GRF53_8_buffer[!clk]) begin
          $fwrite(f, "Register (53,8) Value: %h\n", GRF53_8_buffer[clk]);
        end
        if (GRF53_9_buffer[clk] != GRF53_9_buffer[!clk]) begin
          $fwrite(f, "Register (53,9) Value: %h\n", GRF53_9_buffer[clk]);
        end
        if (GRF53_10_buffer[clk] != GRF53_10_buffer[!clk]) begin
          $fwrite(f, "Register (53,10) Value: %h\n", GRF53_10_buffer[clk]);
        end
        if (GRF53_11_buffer[clk] != GRF53_11_buffer[!clk]) begin
          $fwrite(f, "Register (53,11) Value: %h\n", GRF53_11_buffer[clk]);
        end
        if (GRF53_12_buffer[clk] != GRF53_12_buffer[!clk]) begin
          $fwrite(f, "Register (53,12) Value: %h\n", GRF53_12_buffer[clk]);
        end
        if (GRF53_13_buffer[clk] != GRF53_13_buffer[!clk]) begin
          $fwrite(f, "Register (53,13) Value: %h\n", GRF53_13_buffer[clk]);
        end
        if (GRF53_14_buffer[clk] != GRF53_14_buffer[!clk]) begin
          $fwrite(f, "Register (53,14) Value: %h\n", GRF53_14_buffer[clk]);
        end
        if (GRF53_15_buffer[clk] != GRF53_15_buffer[!clk]) begin
          $fwrite(f, "Register (53,15) Value: %h\n", GRF53_15_buffer[clk]);
        end
        if (GRF53_16_buffer[clk] != GRF53_16_buffer[!clk]) begin
          $fwrite(f, "Register (53,16) Value: %h\n", GRF53_16_buffer[clk]);
        end
        if (GRF53_17_buffer[clk] != GRF53_17_buffer[!clk]) begin
          $fwrite(f, "Register (53,17) Value: %h\n", GRF53_17_buffer[clk]);
        end
        if (GRF53_18_buffer[clk] != GRF53_18_buffer[!clk]) begin
          $fwrite(f, "Register (53,18) Value: %h\n", GRF53_18_buffer[clk]);
        end
        if (GRF53_19_buffer[clk] != GRF53_19_buffer[!clk]) begin
          $fwrite(f, "Register (53,19) Value: %h\n", GRF53_19_buffer[clk]);
        end
        if (GRF53_20_buffer[clk] != GRF53_20_buffer[!clk]) begin
          $fwrite(f, "Register (53,20) Value: %h\n", GRF53_20_buffer[clk]);
        end
        if (GRF53_21_buffer[clk] != GRF53_21_buffer[!clk]) begin
          $fwrite(f, "Register (53,21) Value: %h\n", GRF53_21_buffer[clk]);
        end
        if (GRF53_22_buffer[clk] != GRF53_22_buffer[!clk]) begin
          $fwrite(f, "Register (53,22) Value: %h\n", GRF53_22_buffer[clk]);
        end
        if (GRF53_23_buffer[clk] != GRF53_23_buffer[!clk]) begin
          $fwrite(f, "Register (53,23) Value: %h\n", GRF53_23_buffer[clk]);
        end
        if (GRF53_24_buffer[clk] != GRF53_24_buffer[!clk]) begin
          $fwrite(f, "Register (53,24) Value: %h\n", GRF53_24_buffer[clk]);
        end
        if (GRF53_25_buffer[clk] != GRF53_25_buffer[!clk]) begin
          $fwrite(f, "Register (53,25) Value: %h\n", GRF53_25_buffer[clk]);
        end
        if (GRF53_26_buffer[clk] != GRF53_26_buffer[!clk]) begin
          $fwrite(f, "Register (53,26) Value: %h\n", GRF53_26_buffer[clk]);
        end
        if (GRF53_27_buffer[clk] != GRF53_27_buffer[!clk]) begin
          $fwrite(f, "Register (53,27) Value: %h\n", GRF53_27_buffer[clk]);
        end
        if (GRF53_28_buffer[clk] != GRF53_28_buffer[!clk]) begin
          $fwrite(f, "Register (53,28) Value: %h\n", GRF53_28_buffer[clk]);
        end
        if (GRF53_29_buffer[clk] != GRF53_29_buffer[!clk]) begin
          $fwrite(f, "Register (53,29) Value: %h\n", GRF53_29_buffer[clk]);
        end
        if (GRF53_30_buffer[clk] != GRF53_30_buffer[!clk]) begin
          $fwrite(f, "Register (53,30) Value: %h\n", GRF53_30_buffer[clk]);
        end
        if (GRF53_31_buffer[clk] != GRF53_31_buffer[!clk]) begin
          $fwrite(f, "Register (53,31) Value: %h\n", GRF53_31_buffer[clk]);
        end
        if (GRF54_0_buffer[clk] != GRF54_0_buffer[!clk]) begin
          $fwrite(f, "Register (54,0) Value: %h\n", GRF54_0_buffer[clk]);
        end
        if (GRF54_1_buffer[clk] != GRF54_1_buffer[!clk]) begin
          $fwrite(f, "Register (54,1) Value: %h\n", GRF54_1_buffer[clk]);
        end
        if (GRF54_2_buffer[clk] != GRF54_2_buffer[!clk]) begin
          $fwrite(f, "Register (54,2) Value: %h\n", GRF54_2_buffer[clk]);
        end
        if (GRF54_3_buffer[clk] != GRF54_3_buffer[!clk]) begin
          $fwrite(f, "Register (54,3) Value: %h\n", GRF54_3_buffer[clk]);
        end
        if (GRF54_4_buffer[clk] != GRF54_4_buffer[!clk]) begin
          $fwrite(f, "Register (54,4) Value: %h\n", GRF54_4_buffer[clk]);
        end
        if (GRF54_5_buffer[clk] != GRF54_5_buffer[!clk]) begin
          $fwrite(f, "Register (54,5) Value: %h\n", GRF54_5_buffer[clk]);
        end
        if (GRF54_6_buffer[clk] != GRF54_6_buffer[!clk]) begin
          $fwrite(f, "Register (54,6) Value: %h\n", GRF54_6_buffer[clk]);
        end
        if (GRF54_7_buffer[clk] != GRF54_7_buffer[!clk]) begin
          $fwrite(f, "Register (54,7) Value: %h\n", GRF54_7_buffer[clk]);
        end
        if (GRF54_8_buffer[clk] != GRF54_8_buffer[!clk]) begin
          $fwrite(f, "Register (54,8) Value: %h\n", GRF54_8_buffer[clk]);
        end
        if (GRF54_9_buffer[clk] != GRF54_9_buffer[!clk]) begin
          $fwrite(f, "Register (54,9) Value: %h\n", GRF54_9_buffer[clk]);
        end
        if (GRF54_10_buffer[clk] != GRF54_10_buffer[!clk]) begin
          $fwrite(f, "Register (54,10) Value: %h\n", GRF54_10_buffer[clk]);
        end
        if (GRF54_11_buffer[clk] != GRF54_11_buffer[!clk]) begin
          $fwrite(f, "Register (54,11) Value: %h\n", GRF54_11_buffer[clk]);
        end
        if (GRF54_12_buffer[clk] != GRF54_12_buffer[!clk]) begin
          $fwrite(f, "Register (54,12) Value: %h\n", GRF54_12_buffer[clk]);
        end
        if (GRF54_13_buffer[clk] != GRF54_13_buffer[!clk]) begin
          $fwrite(f, "Register (54,13) Value: %h\n", GRF54_13_buffer[clk]);
        end
        if (GRF54_14_buffer[clk] != GRF54_14_buffer[!clk]) begin
          $fwrite(f, "Register (54,14) Value: %h\n", GRF54_14_buffer[clk]);
        end
        if (GRF54_15_buffer[clk] != GRF54_15_buffer[!clk]) begin
          $fwrite(f, "Register (54,15) Value: %h\n", GRF54_15_buffer[clk]);
        end
        if (GRF54_16_buffer[clk] != GRF54_16_buffer[!clk]) begin
          $fwrite(f, "Register (54,16) Value: %h\n", GRF54_16_buffer[clk]);
        end
        if (GRF54_17_buffer[clk] != GRF54_17_buffer[!clk]) begin
          $fwrite(f, "Register (54,17) Value: %h\n", GRF54_17_buffer[clk]);
        end
        if (GRF54_18_buffer[clk] != GRF54_18_buffer[!clk]) begin
          $fwrite(f, "Register (54,18) Value: %h\n", GRF54_18_buffer[clk]);
        end
        if (GRF54_19_buffer[clk] != GRF54_19_buffer[!clk]) begin
          $fwrite(f, "Register (54,19) Value: %h\n", GRF54_19_buffer[clk]);
        end
        if (GRF54_20_buffer[clk] != GRF54_20_buffer[!clk]) begin
          $fwrite(f, "Register (54,20) Value: %h\n", GRF54_20_buffer[clk]);
        end
        if (GRF54_21_buffer[clk] != GRF54_21_buffer[!clk]) begin
          $fwrite(f, "Register (54,21) Value: %h\n", GRF54_21_buffer[clk]);
        end
        if (GRF54_22_buffer[clk] != GRF54_22_buffer[!clk]) begin
          $fwrite(f, "Register (54,22) Value: %h\n", GRF54_22_buffer[clk]);
        end
        if (GRF54_23_buffer[clk] != GRF54_23_buffer[!clk]) begin
          $fwrite(f, "Register (54,23) Value: %h\n", GRF54_23_buffer[clk]);
        end
        if (GRF54_24_buffer[clk] != GRF54_24_buffer[!clk]) begin
          $fwrite(f, "Register (54,24) Value: %h\n", GRF54_24_buffer[clk]);
        end
        if (GRF54_25_buffer[clk] != GRF54_25_buffer[!clk]) begin
          $fwrite(f, "Register (54,25) Value: %h\n", GRF54_25_buffer[clk]);
        end
        if (GRF54_26_buffer[clk] != GRF54_26_buffer[!clk]) begin
          $fwrite(f, "Register (54,26) Value: %h\n", GRF54_26_buffer[clk]);
        end
        if (GRF54_27_buffer[clk] != GRF54_27_buffer[!clk]) begin
          $fwrite(f, "Register (54,27) Value: %h\n", GRF54_27_buffer[clk]);
        end
        if (GRF54_28_buffer[clk] != GRF54_28_buffer[!clk]) begin
          $fwrite(f, "Register (54,28) Value: %h\n", GRF54_28_buffer[clk]);
        end
        if (GRF54_29_buffer[clk] != GRF54_29_buffer[!clk]) begin
          $fwrite(f, "Register (54,29) Value: %h\n", GRF54_29_buffer[clk]);
        end
        if (GRF54_30_buffer[clk] != GRF54_30_buffer[!clk]) begin
          $fwrite(f, "Register (54,30) Value: %h\n", GRF54_30_buffer[clk]);
        end
        if (GRF54_31_buffer[clk] != GRF54_31_buffer[!clk]) begin
          $fwrite(f, "Register (54,31) Value: %h\n", GRF54_31_buffer[clk]);
        end
        if (GRF55_0_buffer[clk] != GRF55_0_buffer[!clk]) begin
          $fwrite(f, "Register (55,0) Value: %h\n", GRF55_0_buffer[clk]);
        end
        if (GRF55_1_buffer[clk] != GRF55_1_buffer[!clk]) begin
          $fwrite(f, "Register (55,1) Value: %h\n", GRF55_1_buffer[clk]);
        end
        if (GRF55_2_buffer[clk] != GRF55_2_buffer[!clk]) begin
          $fwrite(f, "Register (55,2) Value: %h\n", GRF55_2_buffer[clk]);
        end
        if (GRF55_3_buffer[clk] != GRF55_3_buffer[!clk]) begin
          $fwrite(f, "Register (55,3) Value: %h\n", GRF55_3_buffer[clk]);
        end
        if (GRF55_4_buffer[clk] != GRF55_4_buffer[!clk]) begin
          $fwrite(f, "Register (55,4) Value: %h\n", GRF55_4_buffer[clk]);
        end
        if (GRF55_5_buffer[clk] != GRF55_5_buffer[!clk]) begin
          $fwrite(f, "Register (55,5) Value: %h\n", GRF55_5_buffer[clk]);
        end
        if (GRF55_6_buffer[clk] != GRF55_6_buffer[!clk]) begin
          $fwrite(f, "Register (55,6) Value: %h\n", GRF55_6_buffer[clk]);
        end
        if (GRF55_7_buffer[clk] != GRF55_7_buffer[!clk]) begin
          $fwrite(f, "Register (55,7) Value: %h\n", GRF55_7_buffer[clk]);
        end
        if (GRF55_8_buffer[clk] != GRF55_8_buffer[!clk]) begin
          $fwrite(f, "Register (55,8) Value: %h\n", GRF55_8_buffer[clk]);
        end
        if (GRF55_9_buffer[clk] != GRF55_9_buffer[!clk]) begin
          $fwrite(f, "Register (55,9) Value: %h\n", GRF55_9_buffer[clk]);
        end
        if (GRF55_10_buffer[clk] != GRF55_10_buffer[!clk]) begin
          $fwrite(f, "Register (55,10) Value: %h\n", GRF55_10_buffer[clk]);
        end
        if (GRF55_11_buffer[clk] != GRF55_11_buffer[!clk]) begin
          $fwrite(f, "Register (55,11) Value: %h\n", GRF55_11_buffer[clk]);
        end
        if (GRF55_12_buffer[clk] != GRF55_12_buffer[!clk]) begin
          $fwrite(f, "Register (55,12) Value: %h\n", GRF55_12_buffer[clk]);
        end
        if (GRF55_13_buffer[clk] != GRF55_13_buffer[!clk]) begin
          $fwrite(f, "Register (55,13) Value: %h\n", GRF55_13_buffer[clk]);
        end
        if (GRF55_14_buffer[clk] != GRF55_14_buffer[!clk]) begin
          $fwrite(f, "Register (55,14) Value: %h\n", GRF55_14_buffer[clk]);
        end
        if (GRF55_15_buffer[clk] != GRF55_15_buffer[!clk]) begin
          $fwrite(f, "Register (55,15) Value: %h\n", GRF55_15_buffer[clk]);
        end
        if (GRF55_16_buffer[clk] != GRF55_16_buffer[!clk]) begin
          $fwrite(f, "Register (55,16) Value: %h\n", GRF55_16_buffer[clk]);
        end
        if (GRF55_17_buffer[clk] != GRF55_17_buffer[!clk]) begin
          $fwrite(f, "Register (55,17) Value: %h\n", GRF55_17_buffer[clk]);
        end
        if (GRF55_18_buffer[clk] != GRF55_18_buffer[!clk]) begin
          $fwrite(f, "Register (55,18) Value: %h\n", GRF55_18_buffer[clk]);
        end
        if (GRF55_19_buffer[clk] != GRF55_19_buffer[!clk]) begin
          $fwrite(f, "Register (55,19) Value: %h\n", GRF55_19_buffer[clk]);
        end
        if (GRF55_20_buffer[clk] != GRF55_20_buffer[!clk]) begin
          $fwrite(f, "Register (55,20) Value: %h\n", GRF55_20_buffer[clk]);
        end
        if (GRF55_21_buffer[clk] != GRF55_21_buffer[!clk]) begin
          $fwrite(f, "Register (55,21) Value: %h\n", GRF55_21_buffer[clk]);
        end
        if (GRF55_22_buffer[clk] != GRF55_22_buffer[!clk]) begin
          $fwrite(f, "Register (55,22) Value: %h\n", GRF55_22_buffer[clk]);
        end
        if (GRF55_23_buffer[clk] != GRF55_23_buffer[!clk]) begin
          $fwrite(f, "Register (55,23) Value: %h\n", GRF55_23_buffer[clk]);
        end
        if (GRF55_24_buffer[clk] != GRF55_24_buffer[!clk]) begin
          $fwrite(f, "Register (55,24) Value: %h\n", GRF55_24_buffer[clk]);
        end
        if (GRF55_25_buffer[clk] != GRF55_25_buffer[!clk]) begin
          $fwrite(f, "Register (55,25) Value: %h\n", GRF55_25_buffer[clk]);
        end
        if (GRF55_26_buffer[clk] != GRF55_26_buffer[!clk]) begin
          $fwrite(f, "Register (55,26) Value: %h\n", GRF55_26_buffer[clk]);
        end
        if (GRF55_27_buffer[clk] != GRF55_27_buffer[!clk]) begin
          $fwrite(f, "Register (55,27) Value: %h\n", GRF55_27_buffer[clk]);
        end
        if (GRF55_28_buffer[clk] != GRF55_28_buffer[!clk]) begin
          $fwrite(f, "Register (55,28) Value: %h\n", GRF55_28_buffer[clk]);
        end
        if (GRF55_29_buffer[clk] != GRF55_29_buffer[!clk]) begin
          $fwrite(f, "Register (55,29) Value: %h\n", GRF55_29_buffer[clk]);
        end
        if (GRF55_30_buffer[clk] != GRF55_30_buffer[!clk]) begin
          $fwrite(f, "Register (55,30) Value: %h\n", GRF55_30_buffer[clk]);
        end
        if (GRF55_31_buffer[clk] != GRF55_31_buffer[!clk]) begin
          $fwrite(f, "Register (55,31) Value: %h\n", GRF55_31_buffer[clk]);
        end
        if (GRF56_0_buffer[clk] != GRF56_0_buffer[!clk]) begin
          $fwrite(f, "Register (56,0) Value: %h\n", GRF56_0_buffer[clk]);
        end
        if (GRF56_1_buffer[clk] != GRF56_1_buffer[!clk]) begin
          $fwrite(f, "Register (56,1) Value: %h\n", GRF56_1_buffer[clk]);
        end
        if (GRF56_2_buffer[clk] != GRF56_2_buffer[!clk]) begin
          $fwrite(f, "Register (56,2) Value: %h\n", GRF56_2_buffer[clk]);
        end
        if (GRF56_3_buffer[clk] != GRF56_3_buffer[!clk]) begin
          $fwrite(f, "Register (56,3) Value: %h\n", GRF56_3_buffer[clk]);
        end
        if (GRF56_4_buffer[clk] != GRF56_4_buffer[!clk]) begin
          $fwrite(f, "Register (56,4) Value: %h\n", GRF56_4_buffer[clk]);
        end
        if (GRF56_5_buffer[clk] != GRF56_5_buffer[!clk]) begin
          $fwrite(f, "Register (56,5) Value: %h\n", GRF56_5_buffer[clk]);
        end
        if (GRF56_6_buffer[clk] != GRF56_6_buffer[!clk]) begin
          $fwrite(f, "Register (56,6) Value: %h\n", GRF56_6_buffer[clk]);
        end
        if (GRF56_7_buffer[clk] != GRF56_7_buffer[!clk]) begin
          $fwrite(f, "Register (56,7) Value: %h\n", GRF56_7_buffer[clk]);
        end
        if (GRF56_8_buffer[clk] != GRF56_8_buffer[!clk]) begin
          $fwrite(f, "Register (56,8) Value: %h\n", GRF56_8_buffer[clk]);
        end
        if (GRF56_9_buffer[clk] != GRF56_9_buffer[!clk]) begin
          $fwrite(f, "Register (56,9) Value: %h\n", GRF56_9_buffer[clk]);
        end
        if (GRF56_10_buffer[clk] != GRF56_10_buffer[!clk]) begin
          $fwrite(f, "Register (56,10) Value: %h\n", GRF56_10_buffer[clk]);
        end
        if (GRF56_11_buffer[clk] != GRF56_11_buffer[!clk]) begin
          $fwrite(f, "Register (56,11) Value: %h\n", GRF56_11_buffer[clk]);
        end
        if (GRF56_12_buffer[clk] != GRF56_12_buffer[!clk]) begin
          $fwrite(f, "Register (56,12) Value: %h\n", GRF56_12_buffer[clk]);
        end
        if (GRF56_13_buffer[clk] != GRF56_13_buffer[!clk]) begin
          $fwrite(f, "Register (56,13) Value: %h\n", GRF56_13_buffer[clk]);
        end
        if (GRF56_14_buffer[clk] != GRF56_14_buffer[!clk]) begin
          $fwrite(f, "Register (56,14) Value: %h\n", GRF56_14_buffer[clk]);
        end
        if (GRF56_15_buffer[clk] != GRF56_15_buffer[!clk]) begin
          $fwrite(f, "Register (56,15) Value: %h\n", GRF56_15_buffer[clk]);
        end
        if (GRF56_16_buffer[clk] != GRF56_16_buffer[!clk]) begin
          $fwrite(f, "Register (56,16) Value: %h\n", GRF56_16_buffer[clk]);
        end
        if (GRF56_17_buffer[clk] != GRF56_17_buffer[!clk]) begin
          $fwrite(f, "Register (56,17) Value: %h\n", GRF56_17_buffer[clk]);
        end
        if (GRF56_18_buffer[clk] != GRF56_18_buffer[!clk]) begin
          $fwrite(f, "Register (56,18) Value: %h\n", GRF56_18_buffer[clk]);
        end
        if (GRF56_19_buffer[clk] != GRF56_19_buffer[!clk]) begin
          $fwrite(f, "Register (56,19) Value: %h\n", GRF56_19_buffer[clk]);
        end
        if (GRF56_20_buffer[clk] != GRF56_20_buffer[!clk]) begin
          $fwrite(f, "Register (56,20) Value: %h\n", GRF56_20_buffer[clk]);
        end
        if (GRF56_21_buffer[clk] != GRF56_21_buffer[!clk]) begin
          $fwrite(f, "Register (56,21) Value: %h\n", GRF56_21_buffer[clk]);
        end
        if (GRF56_22_buffer[clk] != GRF56_22_buffer[!clk]) begin
          $fwrite(f, "Register (56,22) Value: %h\n", GRF56_22_buffer[clk]);
        end
        if (GRF56_23_buffer[clk] != GRF56_23_buffer[!clk]) begin
          $fwrite(f, "Register (56,23) Value: %h\n", GRF56_23_buffer[clk]);
        end
        if (GRF56_24_buffer[clk] != GRF56_24_buffer[!clk]) begin
          $fwrite(f, "Register (56,24) Value: %h\n", GRF56_24_buffer[clk]);
        end
        if (GRF56_25_buffer[clk] != GRF56_25_buffer[!clk]) begin
          $fwrite(f, "Register (56,25) Value: %h\n", GRF56_25_buffer[clk]);
        end
        if (GRF56_26_buffer[clk] != GRF56_26_buffer[!clk]) begin
          $fwrite(f, "Register (56,26) Value: %h\n", GRF56_26_buffer[clk]);
        end
        if (GRF56_27_buffer[clk] != GRF56_27_buffer[!clk]) begin
          $fwrite(f, "Register (56,27) Value: %h\n", GRF56_27_buffer[clk]);
        end
        if (GRF56_28_buffer[clk] != GRF56_28_buffer[!clk]) begin
          $fwrite(f, "Register (56,28) Value: %h\n", GRF56_28_buffer[clk]);
        end
        if (GRF56_29_buffer[clk] != GRF56_29_buffer[!clk]) begin
          $fwrite(f, "Register (56,29) Value: %h\n", GRF56_29_buffer[clk]);
        end
        if (GRF56_30_buffer[clk] != GRF56_30_buffer[!clk]) begin
          $fwrite(f, "Register (56,30) Value: %h\n", GRF56_30_buffer[clk]);
        end
        if (GRF56_31_buffer[clk] != GRF56_31_buffer[!clk]) begin
          $fwrite(f, "Register (56,31) Value: %h\n", GRF56_31_buffer[clk]);
        end
        if (GRF57_0_buffer[clk] != GRF57_0_buffer[!clk]) begin
          $fwrite(f, "Register (57,0) Value: %h\n", GRF57_0_buffer[clk]);
        end
        if (GRF57_1_buffer[clk] != GRF57_1_buffer[!clk]) begin
          $fwrite(f, "Register (57,1) Value: %h\n", GRF57_1_buffer[clk]);
        end
        if (GRF57_2_buffer[clk] != GRF57_2_buffer[!clk]) begin
          $fwrite(f, "Register (57,2) Value: %h\n", GRF57_2_buffer[clk]);
        end
        if (GRF57_3_buffer[clk] != GRF57_3_buffer[!clk]) begin
          $fwrite(f, "Register (57,3) Value: %h\n", GRF57_3_buffer[clk]);
        end
        if (GRF57_4_buffer[clk] != GRF57_4_buffer[!clk]) begin
          $fwrite(f, "Register (57,4) Value: %h\n", GRF57_4_buffer[clk]);
        end
        if (GRF57_5_buffer[clk] != GRF57_5_buffer[!clk]) begin
          $fwrite(f, "Register (57,5) Value: %h\n", GRF57_5_buffer[clk]);
        end
        if (GRF57_6_buffer[clk] != GRF57_6_buffer[!clk]) begin
          $fwrite(f, "Register (57,6) Value: %h\n", GRF57_6_buffer[clk]);
        end
        if (GRF57_7_buffer[clk] != GRF57_7_buffer[!clk]) begin
          $fwrite(f, "Register (57,7) Value: %h\n", GRF57_7_buffer[clk]);
        end
        if (GRF57_8_buffer[clk] != GRF57_8_buffer[!clk]) begin
          $fwrite(f, "Register (57,8) Value: %h\n", GRF57_8_buffer[clk]);
        end
        if (GRF57_9_buffer[clk] != GRF57_9_buffer[!clk]) begin
          $fwrite(f, "Register (57,9) Value: %h\n", GRF57_9_buffer[clk]);
        end
        if (GRF57_10_buffer[clk] != GRF57_10_buffer[!clk]) begin
          $fwrite(f, "Register (57,10) Value: %h\n", GRF57_10_buffer[clk]);
        end
        if (GRF57_11_buffer[clk] != GRF57_11_buffer[!clk]) begin
          $fwrite(f, "Register (57,11) Value: %h\n", GRF57_11_buffer[clk]);
        end
        if (GRF57_12_buffer[clk] != GRF57_12_buffer[!clk]) begin
          $fwrite(f, "Register (57,12) Value: %h\n", GRF57_12_buffer[clk]);
        end
        if (GRF57_13_buffer[clk] != GRF57_13_buffer[!clk]) begin
          $fwrite(f, "Register (57,13) Value: %h\n", GRF57_13_buffer[clk]);
        end
        if (GRF57_14_buffer[clk] != GRF57_14_buffer[!clk]) begin
          $fwrite(f, "Register (57,14) Value: %h\n", GRF57_14_buffer[clk]);
        end
        if (GRF57_15_buffer[clk] != GRF57_15_buffer[!clk]) begin
          $fwrite(f, "Register (57,15) Value: %h\n", GRF57_15_buffer[clk]);
        end
        if (GRF57_16_buffer[clk] != GRF57_16_buffer[!clk]) begin
          $fwrite(f, "Register (57,16) Value: %h\n", GRF57_16_buffer[clk]);
        end
        if (GRF57_17_buffer[clk] != GRF57_17_buffer[!clk]) begin
          $fwrite(f, "Register (57,17) Value: %h\n", GRF57_17_buffer[clk]);
        end
        if (GRF57_18_buffer[clk] != GRF57_18_buffer[!clk]) begin
          $fwrite(f, "Register (57,18) Value: %h\n", GRF57_18_buffer[clk]);
        end
        if (GRF57_19_buffer[clk] != GRF57_19_buffer[!clk]) begin
          $fwrite(f, "Register (57,19) Value: %h\n", GRF57_19_buffer[clk]);
        end
        if (GRF57_20_buffer[clk] != GRF57_20_buffer[!clk]) begin
          $fwrite(f, "Register (57,20) Value: %h\n", GRF57_20_buffer[clk]);
        end
        if (GRF57_21_buffer[clk] != GRF57_21_buffer[!clk]) begin
          $fwrite(f, "Register (57,21) Value: %h\n", GRF57_21_buffer[clk]);
        end
        if (GRF57_22_buffer[clk] != GRF57_22_buffer[!clk]) begin
          $fwrite(f, "Register (57,22) Value: %h\n", GRF57_22_buffer[clk]);
        end
        if (GRF57_23_buffer[clk] != GRF57_23_buffer[!clk]) begin
          $fwrite(f, "Register (57,23) Value: %h\n", GRF57_23_buffer[clk]);
        end
        if (GRF57_24_buffer[clk] != GRF57_24_buffer[!clk]) begin
          $fwrite(f, "Register (57,24) Value: %h\n", GRF57_24_buffer[clk]);
        end
        if (GRF57_25_buffer[clk] != GRF57_25_buffer[!clk]) begin
          $fwrite(f, "Register (57,25) Value: %h\n", GRF57_25_buffer[clk]);
        end
        if (GRF57_26_buffer[clk] != GRF57_26_buffer[!clk]) begin
          $fwrite(f, "Register (57,26) Value: %h\n", GRF57_26_buffer[clk]);
        end
        if (GRF57_27_buffer[clk] != GRF57_27_buffer[!clk]) begin
          $fwrite(f, "Register (57,27) Value: %h\n", GRF57_27_buffer[clk]);
        end
        if (GRF57_28_buffer[clk] != GRF57_28_buffer[!clk]) begin
          $fwrite(f, "Register (57,28) Value: %h\n", GRF57_28_buffer[clk]);
        end
        if (GRF57_29_buffer[clk] != GRF57_29_buffer[!clk]) begin
          $fwrite(f, "Register (57,29) Value: %h\n", GRF57_29_buffer[clk]);
        end
        if (GRF57_30_buffer[clk] != GRF57_30_buffer[!clk]) begin
          $fwrite(f, "Register (57,30) Value: %h\n", GRF57_30_buffer[clk]);
        end
        if (GRF57_31_buffer[clk] != GRF57_31_buffer[!clk]) begin
          $fwrite(f, "Register (57,31) Value: %h\n", GRF57_31_buffer[clk]);
        end
        if (GRF58_0_buffer[clk] != GRF58_0_buffer[!clk]) begin
          $fwrite(f, "Register (58,0) Value: %h\n", GRF58_0_buffer[clk]);
        end
        if (GRF58_1_buffer[clk] != GRF58_1_buffer[!clk]) begin
          $fwrite(f, "Register (58,1) Value: %h\n", GRF58_1_buffer[clk]);
        end
        if (GRF58_2_buffer[clk] != GRF58_2_buffer[!clk]) begin
          $fwrite(f, "Register (58,2) Value: %h\n", GRF58_2_buffer[clk]);
        end
        if (GRF58_3_buffer[clk] != GRF58_3_buffer[!clk]) begin
          $fwrite(f, "Register (58,3) Value: %h\n", GRF58_3_buffer[clk]);
        end
        if (GRF58_4_buffer[clk] != GRF58_4_buffer[!clk]) begin
          $fwrite(f, "Register (58,4) Value: %h\n", GRF58_4_buffer[clk]);
        end
        if (GRF58_5_buffer[clk] != GRF58_5_buffer[!clk]) begin
          $fwrite(f, "Register (58,5) Value: %h\n", GRF58_5_buffer[clk]);
        end
        if (GRF58_6_buffer[clk] != GRF58_6_buffer[!clk]) begin
          $fwrite(f, "Register (58,6) Value: %h\n", GRF58_6_buffer[clk]);
        end
        if (GRF58_7_buffer[clk] != GRF58_7_buffer[!clk]) begin
          $fwrite(f, "Register (58,7) Value: %h\n", GRF58_7_buffer[clk]);
        end
        if (GRF58_8_buffer[clk] != GRF58_8_buffer[!clk]) begin
          $fwrite(f, "Register (58,8) Value: %h\n", GRF58_8_buffer[clk]);
        end
        if (GRF58_9_buffer[clk] != GRF58_9_buffer[!clk]) begin
          $fwrite(f, "Register (58,9) Value: %h\n", GRF58_9_buffer[clk]);
        end
        if (GRF58_10_buffer[clk] != GRF58_10_buffer[!clk]) begin
          $fwrite(f, "Register (58,10) Value: %h\n", GRF58_10_buffer[clk]);
        end
        if (GRF58_11_buffer[clk] != GRF58_11_buffer[!clk]) begin
          $fwrite(f, "Register (58,11) Value: %h\n", GRF58_11_buffer[clk]);
        end
        if (GRF58_12_buffer[clk] != GRF58_12_buffer[!clk]) begin
          $fwrite(f, "Register (58,12) Value: %h\n", GRF58_12_buffer[clk]);
        end
        if (GRF58_13_buffer[clk] != GRF58_13_buffer[!clk]) begin
          $fwrite(f, "Register (58,13) Value: %h\n", GRF58_13_buffer[clk]);
        end
        if (GRF58_14_buffer[clk] != GRF58_14_buffer[!clk]) begin
          $fwrite(f, "Register (58,14) Value: %h\n", GRF58_14_buffer[clk]);
        end
        if (GRF58_15_buffer[clk] != GRF58_15_buffer[!clk]) begin
          $fwrite(f, "Register (58,15) Value: %h\n", GRF58_15_buffer[clk]);
        end
        if (GRF58_16_buffer[clk] != GRF58_16_buffer[!clk]) begin
          $fwrite(f, "Register (58,16) Value: %h\n", GRF58_16_buffer[clk]);
        end
        if (GRF58_17_buffer[clk] != GRF58_17_buffer[!clk]) begin
          $fwrite(f, "Register (58,17) Value: %h\n", GRF58_17_buffer[clk]);
        end
        if (GRF58_18_buffer[clk] != GRF58_18_buffer[!clk]) begin
          $fwrite(f, "Register (58,18) Value: %h\n", GRF58_18_buffer[clk]);
        end
        if (GRF58_19_buffer[clk] != GRF58_19_buffer[!clk]) begin
          $fwrite(f, "Register (58,19) Value: %h\n", GRF58_19_buffer[clk]);
        end
        if (GRF58_20_buffer[clk] != GRF58_20_buffer[!clk]) begin
          $fwrite(f, "Register (58,20) Value: %h\n", GRF58_20_buffer[clk]);
        end
        if (GRF58_21_buffer[clk] != GRF58_21_buffer[!clk]) begin
          $fwrite(f, "Register (58,21) Value: %h\n", GRF58_21_buffer[clk]);
        end
        if (GRF58_22_buffer[clk] != GRF58_22_buffer[!clk]) begin
          $fwrite(f, "Register (58,22) Value: %h\n", GRF58_22_buffer[clk]);
        end
        if (GRF58_23_buffer[clk] != GRF58_23_buffer[!clk]) begin
          $fwrite(f, "Register (58,23) Value: %h\n", GRF58_23_buffer[clk]);
        end
        if (GRF58_24_buffer[clk] != GRF58_24_buffer[!clk]) begin
          $fwrite(f, "Register (58,24) Value: %h\n", GRF58_24_buffer[clk]);
        end
        if (GRF58_25_buffer[clk] != GRF58_25_buffer[!clk]) begin
          $fwrite(f, "Register (58,25) Value: %h\n", GRF58_25_buffer[clk]);
        end
        if (GRF58_26_buffer[clk] != GRF58_26_buffer[!clk]) begin
          $fwrite(f, "Register (58,26) Value: %h\n", GRF58_26_buffer[clk]);
        end
        if (GRF58_27_buffer[clk] != GRF58_27_buffer[!clk]) begin
          $fwrite(f, "Register (58,27) Value: %h\n", GRF58_27_buffer[clk]);
        end
        if (GRF58_28_buffer[clk] != GRF58_28_buffer[!clk]) begin
          $fwrite(f, "Register (58,28) Value: %h\n", GRF58_28_buffer[clk]);
        end
        if (GRF58_29_buffer[clk] != GRF58_29_buffer[!clk]) begin
          $fwrite(f, "Register (58,29) Value: %h\n", GRF58_29_buffer[clk]);
        end
        if (GRF58_30_buffer[clk] != GRF58_30_buffer[!clk]) begin
          $fwrite(f, "Register (58,30) Value: %h\n", GRF58_30_buffer[clk]);
        end
        if (GRF58_31_buffer[clk] != GRF58_31_buffer[!clk]) begin
          $fwrite(f, "Register (58,31) Value: %h\n", GRF58_31_buffer[clk]);
        end
        if (GRF59_0_buffer[clk] != GRF59_0_buffer[!clk]) begin
          $fwrite(f, "Register (59,0) Value: %h\n", GRF59_0_buffer[clk]);
        end
        if (GRF59_1_buffer[clk] != GRF59_1_buffer[!clk]) begin
          $fwrite(f, "Register (59,1) Value: %h\n", GRF59_1_buffer[clk]);
        end
        if (GRF59_2_buffer[clk] != GRF59_2_buffer[!clk]) begin
          $fwrite(f, "Register (59,2) Value: %h\n", GRF59_2_buffer[clk]);
        end
        if (GRF59_3_buffer[clk] != GRF59_3_buffer[!clk]) begin
          $fwrite(f, "Register (59,3) Value: %h\n", GRF59_3_buffer[clk]);
        end
        if (GRF59_4_buffer[clk] != GRF59_4_buffer[!clk]) begin
          $fwrite(f, "Register (59,4) Value: %h\n", GRF59_4_buffer[clk]);
        end
        if (GRF59_5_buffer[clk] != GRF59_5_buffer[!clk]) begin
          $fwrite(f, "Register (59,5) Value: %h\n", GRF59_5_buffer[clk]);
        end
        if (GRF59_6_buffer[clk] != GRF59_6_buffer[!clk]) begin
          $fwrite(f, "Register (59,6) Value: %h\n", GRF59_6_buffer[clk]);
        end
        if (GRF59_7_buffer[clk] != GRF59_7_buffer[!clk]) begin
          $fwrite(f, "Register (59,7) Value: %h\n", GRF59_7_buffer[clk]);
        end
        if (GRF59_8_buffer[clk] != GRF59_8_buffer[!clk]) begin
          $fwrite(f, "Register (59,8) Value: %h\n", GRF59_8_buffer[clk]);
        end
        if (GRF59_9_buffer[clk] != GRF59_9_buffer[!clk]) begin
          $fwrite(f, "Register (59,9) Value: %h\n", GRF59_9_buffer[clk]);
        end
        if (GRF59_10_buffer[clk] != GRF59_10_buffer[!clk]) begin
          $fwrite(f, "Register (59,10) Value: %h\n", GRF59_10_buffer[clk]);
        end
        if (GRF59_11_buffer[clk] != GRF59_11_buffer[!clk]) begin
          $fwrite(f, "Register (59,11) Value: %h\n", GRF59_11_buffer[clk]);
        end
        if (GRF59_12_buffer[clk] != GRF59_12_buffer[!clk]) begin
          $fwrite(f, "Register (59,12) Value: %h\n", GRF59_12_buffer[clk]);
        end
        if (GRF59_13_buffer[clk] != GRF59_13_buffer[!clk]) begin
          $fwrite(f, "Register (59,13) Value: %h\n", GRF59_13_buffer[clk]);
        end
        if (GRF59_14_buffer[clk] != GRF59_14_buffer[!clk]) begin
          $fwrite(f, "Register (59,14) Value: %h\n", GRF59_14_buffer[clk]);
        end
        if (GRF59_15_buffer[clk] != GRF59_15_buffer[!clk]) begin
          $fwrite(f, "Register (59,15) Value: %h\n", GRF59_15_buffer[clk]);
        end
        if (GRF59_16_buffer[clk] != GRF59_16_buffer[!clk]) begin
          $fwrite(f, "Register (59,16) Value: %h\n", GRF59_16_buffer[clk]);
        end
        if (GRF59_17_buffer[clk] != GRF59_17_buffer[!clk]) begin
          $fwrite(f, "Register (59,17) Value: %h\n", GRF59_17_buffer[clk]);
        end
        if (GRF59_18_buffer[clk] != GRF59_18_buffer[!clk]) begin
          $fwrite(f, "Register (59,18) Value: %h\n", GRF59_18_buffer[clk]);
        end
        if (GRF59_19_buffer[clk] != GRF59_19_buffer[!clk]) begin
          $fwrite(f, "Register (59,19) Value: %h\n", GRF59_19_buffer[clk]);
        end
        if (GRF59_20_buffer[clk] != GRF59_20_buffer[!clk]) begin
          $fwrite(f, "Register (59,20) Value: %h\n", GRF59_20_buffer[clk]);
        end
        if (GRF59_21_buffer[clk] != GRF59_21_buffer[!clk]) begin
          $fwrite(f, "Register (59,21) Value: %h\n", GRF59_21_buffer[clk]);
        end
        if (GRF59_22_buffer[clk] != GRF59_22_buffer[!clk]) begin
          $fwrite(f, "Register (59,22) Value: %h\n", GRF59_22_buffer[clk]);
        end
        if (GRF59_23_buffer[clk] != GRF59_23_buffer[!clk]) begin
          $fwrite(f, "Register (59,23) Value: %h\n", GRF59_23_buffer[clk]);
        end
        if (GRF59_24_buffer[clk] != GRF59_24_buffer[!clk]) begin
          $fwrite(f, "Register (59,24) Value: %h\n", GRF59_24_buffer[clk]);
        end
        if (GRF59_25_buffer[clk] != GRF59_25_buffer[!clk]) begin
          $fwrite(f, "Register (59,25) Value: %h\n", GRF59_25_buffer[clk]);
        end
        if (GRF59_26_buffer[clk] != GRF59_26_buffer[!clk]) begin
          $fwrite(f, "Register (59,26) Value: %h\n", GRF59_26_buffer[clk]);
        end
        if (GRF59_27_buffer[clk] != GRF59_27_buffer[!clk]) begin
          $fwrite(f, "Register (59,27) Value: %h\n", GRF59_27_buffer[clk]);
        end
        if (GRF59_28_buffer[clk] != GRF59_28_buffer[!clk]) begin
          $fwrite(f, "Register (59,28) Value: %h\n", GRF59_28_buffer[clk]);
        end
        if (GRF59_29_buffer[clk] != GRF59_29_buffer[!clk]) begin
          $fwrite(f, "Register (59,29) Value: %h\n", GRF59_29_buffer[clk]);
        end
        if (GRF59_30_buffer[clk] != GRF59_30_buffer[!clk]) begin
          $fwrite(f, "Register (59,30) Value: %h\n", GRF59_30_buffer[clk]);
        end
        if (GRF59_31_buffer[clk] != GRF59_31_buffer[!clk]) begin
          $fwrite(f, "Register (59,31) Value: %h\n", GRF59_31_buffer[clk]);
        end
        if (GRF60_0_buffer[clk] != GRF60_0_buffer[!clk]) begin
          $fwrite(f, "Register (60,0) Value: %h\n", GRF60_0_buffer[clk]);
        end
        if (GRF60_1_buffer[clk] != GRF60_1_buffer[!clk]) begin
          $fwrite(f, "Register (60,1) Value: %h\n", GRF60_1_buffer[clk]);
        end
        if (GRF60_2_buffer[clk] != GRF60_2_buffer[!clk]) begin
          $fwrite(f, "Register (60,2) Value: %h\n", GRF60_2_buffer[clk]);
        end
        if (GRF60_3_buffer[clk] != GRF60_3_buffer[!clk]) begin
          $fwrite(f, "Register (60,3) Value: %h\n", GRF60_3_buffer[clk]);
        end
        if (GRF60_4_buffer[clk] != GRF60_4_buffer[!clk]) begin
          $fwrite(f, "Register (60,4) Value: %h\n", GRF60_4_buffer[clk]);
        end
        if (GRF60_5_buffer[clk] != GRF60_5_buffer[!clk]) begin
          $fwrite(f, "Register (60,5) Value: %h\n", GRF60_5_buffer[clk]);
        end
        if (GRF60_6_buffer[clk] != GRF60_6_buffer[!clk]) begin
          $fwrite(f, "Register (60,6) Value: %h\n", GRF60_6_buffer[clk]);
        end
        if (GRF60_7_buffer[clk] != GRF60_7_buffer[!clk]) begin
          $fwrite(f, "Register (60,7) Value: %h\n", GRF60_7_buffer[clk]);
        end
        if (GRF60_8_buffer[clk] != GRF60_8_buffer[!clk]) begin
          $fwrite(f, "Register (60,8) Value: %h\n", GRF60_8_buffer[clk]);
        end
        if (GRF60_9_buffer[clk] != GRF60_9_buffer[!clk]) begin
          $fwrite(f, "Register (60,9) Value: %h\n", GRF60_9_buffer[clk]);
        end
        if (GRF60_10_buffer[clk] != GRF60_10_buffer[!clk]) begin
          $fwrite(f, "Register (60,10) Value: %h\n", GRF60_10_buffer[clk]);
        end
        if (GRF60_11_buffer[clk] != GRF60_11_buffer[!clk]) begin
          $fwrite(f, "Register (60,11) Value: %h\n", GRF60_11_buffer[clk]);
        end
        if (GRF60_12_buffer[clk] != GRF60_12_buffer[!clk]) begin
          $fwrite(f, "Register (60,12) Value: %h\n", GRF60_12_buffer[clk]);
        end
        if (GRF60_13_buffer[clk] != GRF60_13_buffer[!clk]) begin
          $fwrite(f, "Register (60,13) Value: %h\n", GRF60_13_buffer[clk]);
        end
        if (GRF60_14_buffer[clk] != GRF60_14_buffer[!clk]) begin
          $fwrite(f, "Register (60,14) Value: %h\n", GRF60_14_buffer[clk]);
        end
        if (GRF60_15_buffer[clk] != GRF60_15_buffer[!clk]) begin
          $fwrite(f, "Register (60,15) Value: %h\n", GRF60_15_buffer[clk]);
        end
        if (GRF60_16_buffer[clk] != GRF60_16_buffer[!clk]) begin
          $fwrite(f, "Register (60,16) Value: %h\n", GRF60_16_buffer[clk]);
        end
        if (GRF60_17_buffer[clk] != GRF60_17_buffer[!clk]) begin
          $fwrite(f, "Register (60,17) Value: %h\n", GRF60_17_buffer[clk]);
        end
        if (GRF60_18_buffer[clk] != GRF60_18_buffer[!clk]) begin
          $fwrite(f, "Register (60,18) Value: %h\n", GRF60_18_buffer[clk]);
        end
        if (GRF60_19_buffer[clk] != GRF60_19_buffer[!clk]) begin
          $fwrite(f, "Register (60,19) Value: %h\n", GRF60_19_buffer[clk]);
        end
        if (GRF60_20_buffer[clk] != GRF60_20_buffer[!clk]) begin
          $fwrite(f, "Register (60,20) Value: %h\n", GRF60_20_buffer[clk]);
        end
        if (GRF60_21_buffer[clk] != GRF60_21_buffer[!clk]) begin
          $fwrite(f, "Register (60,21) Value: %h\n", GRF60_21_buffer[clk]);
        end
        if (GRF60_22_buffer[clk] != GRF60_22_buffer[!clk]) begin
          $fwrite(f, "Register (60,22) Value: %h\n", GRF60_22_buffer[clk]);
        end
        if (GRF60_23_buffer[clk] != GRF60_23_buffer[!clk]) begin
          $fwrite(f, "Register (60,23) Value: %h\n", GRF60_23_buffer[clk]);
        end
        if (GRF60_24_buffer[clk] != GRF60_24_buffer[!clk]) begin
          $fwrite(f, "Register (60,24) Value: %h\n", GRF60_24_buffer[clk]);
        end
        if (GRF60_25_buffer[clk] != GRF60_25_buffer[!clk]) begin
          $fwrite(f, "Register (60,25) Value: %h\n", GRF60_25_buffer[clk]);
        end
        if (GRF60_26_buffer[clk] != GRF60_26_buffer[!clk]) begin
          $fwrite(f, "Register (60,26) Value: %h\n", GRF60_26_buffer[clk]);
        end
        if (GRF60_27_buffer[clk] != GRF60_27_buffer[!clk]) begin
          $fwrite(f, "Register (60,27) Value: %h\n", GRF60_27_buffer[clk]);
        end
        if (GRF60_28_buffer[clk] != GRF60_28_buffer[!clk]) begin
          $fwrite(f, "Register (60,28) Value: %h\n", GRF60_28_buffer[clk]);
        end
        if (GRF60_29_buffer[clk] != GRF60_29_buffer[!clk]) begin
          $fwrite(f, "Register (60,29) Value: %h\n", GRF60_29_buffer[clk]);
        end
        if (GRF60_30_buffer[clk] != GRF60_30_buffer[!clk]) begin
          $fwrite(f, "Register (60,30) Value: %h\n", GRF60_30_buffer[clk]);
        end
        if (GRF60_31_buffer[clk] != GRF60_31_buffer[!clk]) begin
          $fwrite(f, "Register (60,31) Value: %h\n", GRF60_31_buffer[clk]);
        end
        if (GRF61_0_buffer[clk] != GRF61_0_buffer[!clk]) begin
          $fwrite(f, "Register (61,0) Value: %h\n", GRF61_0_buffer[clk]);
        end
        if (GRF61_1_buffer[clk] != GRF61_1_buffer[!clk]) begin
          $fwrite(f, "Register (61,1) Value: %h\n", GRF61_1_buffer[clk]);
        end
        if (GRF61_2_buffer[clk] != GRF61_2_buffer[!clk]) begin
          $fwrite(f, "Register (61,2) Value: %h\n", GRF61_2_buffer[clk]);
        end
        if (GRF61_3_buffer[clk] != GRF61_3_buffer[!clk]) begin
          $fwrite(f, "Register (61,3) Value: %h\n", GRF61_3_buffer[clk]);
        end
        if (GRF61_4_buffer[clk] != GRF61_4_buffer[!clk]) begin
          $fwrite(f, "Register (61,4) Value: %h\n", GRF61_4_buffer[clk]);
        end
        if (GRF61_5_buffer[clk] != GRF61_5_buffer[!clk]) begin
          $fwrite(f, "Register (61,5) Value: %h\n", GRF61_5_buffer[clk]);
        end
        if (GRF61_6_buffer[clk] != GRF61_6_buffer[!clk]) begin
          $fwrite(f, "Register (61,6) Value: %h\n", GRF61_6_buffer[clk]);
        end
        if (GRF61_7_buffer[clk] != GRF61_7_buffer[!clk]) begin
          $fwrite(f, "Register (61,7) Value: %h\n", GRF61_7_buffer[clk]);
        end
        if (GRF61_8_buffer[clk] != GRF61_8_buffer[!clk]) begin
          $fwrite(f, "Register (61,8) Value: %h\n", GRF61_8_buffer[clk]);
        end
        if (GRF61_9_buffer[clk] != GRF61_9_buffer[!clk]) begin
          $fwrite(f, "Register (61,9) Value: %h\n", GRF61_9_buffer[clk]);
        end
        if (GRF61_10_buffer[clk] != GRF61_10_buffer[!clk]) begin
          $fwrite(f, "Register (61,10) Value: %h\n", GRF61_10_buffer[clk]);
        end
        if (GRF61_11_buffer[clk] != GRF61_11_buffer[!clk]) begin
          $fwrite(f, "Register (61,11) Value: %h\n", GRF61_11_buffer[clk]);
        end
        if (GRF61_12_buffer[clk] != GRF61_12_buffer[!clk]) begin
          $fwrite(f, "Register (61,12) Value: %h\n", GRF61_12_buffer[clk]);
        end
        if (GRF61_13_buffer[clk] != GRF61_13_buffer[!clk]) begin
          $fwrite(f, "Register (61,13) Value: %h\n", GRF61_13_buffer[clk]);
        end
        if (GRF61_14_buffer[clk] != GRF61_14_buffer[!clk]) begin
          $fwrite(f, "Register (61,14) Value: %h\n", GRF61_14_buffer[clk]);
        end
        if (GRF61_15_buffer[clk] != GRF61_15_buffer[!clk]) begin
          $fwrite(f, "Register (61,15) Value: %h\n", GRF61_15_buffer[clk]);
        end
        if (GRF61_16_buffer[clk] != GRF61_16_buffer[!clk]) begin
          $fwrite(f, "Register (61,16) Value: %h\n", GRF61_16_buffer[clk]);
        end
        if (GRF61_17_buffer[clk] != GRF61_17_buffer[!clk]) begin
          $fwrite(f, "Register (61,17) Value: %h\n", GRF61_17_buffer[clk]);
        end
        if (GRF61_18_buffer[clk] != GRF61_18_buffer[!clk]) begin
          $fwrite(f, "Register (61,18) Value: %h\n", GRF61_18_buffer[clk]);
        end
        if (GRF61_19_buffer[clk] != GRF61_19_buffer[!clk]) begin
          $fwrite(f, "Register (61,19) Value: %h\n", GRF61_19_buffer[clk]);
        end
        if (GRF61_20_buffer[clk] != GRF61_20_buffer[!clk]) begin
          $fwrite(f, "Register (61,20) Value: %h\n", GRF61_20_buffer[clk]);
        end
        if (GRF61_21_buffer[clk] != GRF61_21_buffer[!clk]) begin
          $fwrite(f, "Register (61,21) Value: %h\n", GRF61_21_buffer[clk]);
        end
        if (GRF61_22_buffer[clk] != GRF61_22_buffer[!clk]) begin
          $fwrite(f, "Register (61,22) Value: %h\n", GRF61_22_buffer[clk]);
        end
        if (GRF61_23_buffer[clk] != GRF61_23_buffer[!clk]) begin
          $fwrite(f, "Register (61,23) Value: %h\n", GRF61_23_buffer[clk]);
        end
        if (GRF61_24_buffer[clk] != GRF61_24_buffer[!clk]) begin
          $fwrite(f, "Register (61,24) Value: %h\n", GRF61_24_buffer[clk]);
        end
        if (GRF61_25_buffer[clk] != GRF61_25_buffer[!clk]) begin
          $fwrite(f, "Register (61,25) Value: %h\n", GRF61_25_buffer[clk]);
        end
        if (GRF61_26_buffer[clk] != GRF61_26_buffer[!clk]) begin
          $fwrite(f, "Register (61,26) Value: %h\n", GRF61_26_buffer[clk]);
        end
        if (GRF61_27_buffer[clk] != GRF61_27_buffer[!clk]) begin
          $fwrite(f, "Register (61,27) Value: %h\n", GRF61_27_buffer[clk]);
        end
        if (GRF61_28_buffer[clk] != GRF61_28_buffer[!clk]) begin
          $fwrite(f, "Register (61,28) Value: %h\n", GRF61_28_buffer[clk]);
        end
        if (GRF61_29_buffer[clk] != GRF61_29_buffer[!clk]) begin
          $fwrite(f, "Register (61,29) Value: %h\n", GRF61_29_buffer[clk]);
        end
        if (GRF61_30_buffer[clk] != GRF61_30_buffer[!clk]) begin
          $fwrite(f, "Register (61,30) Value: %h\n", GRF61_30_buffer[clk]);
        end
        if (GRF61_31_buffer[clk] != GRF61_31_buffer[!clk]) begin
          $fwrite(f, "Register (61,31) Value: %h\n", GRF61_31_buffer[clk]);
        end
        if (GRF62_0_buffer[clk] != GRF62_0_buffer[!clk]) begin
          $fwrite(f, "Register (62,0) Value: %h\n", GRF62_0_buffer[clk]);
        end
        if (GRF62_1_buffer[clk] != GRF62_1_buffer[!clk]) begin
          $fwrite(f, "Register (62,1) Value: %h\n", GRF62_1_buffer[clk]);
        end
        if (GRF62_2_buffer[clk] != GRF62_2_buffer[!clk]) begin
          $fwrite(f, "Register (62,2) Value: %h\n", GRF62_2_buffer[clk]);
        end
        if (GRF62_3_buffer[clk] != GRF62_3_buffer[!clk]) begin
          $fwrite(f, "Register (62,3) Value: %h\n", GRF62_3_buffer[clk]);
        end
        if (GRF62_4_buffer[clk] != GRF62_4_buffer[!clk]) begin
          $fwrite(f, "Register (62,4) Value: %h\n", GRF62_4_buffer[clk]);
        end
        if (GRF62_5_buffer[clk] != GRF62_5_buffer[!clk]) begin
          $fwrite(f, "Register (62,5) Value: %h\n", GRF62_5_buffer[clk]);
        end
        if (GRF62_6_buffer[clk] != GRF62_6_buffer[!clk]) begin
          $fwrite(f, "Register (62,6) Value: %h\n", GRF62_6_buffer[clk]);
        end
        if (GRF62_7_buffer[clk] != GRF62_7_buffer[!clk]) begin
          $fwrite(f, "Register (62,7) Value: %h\n", GRF62_7_buffer[clk]);
        end
        if (GRF62_8_buffer[clk] != GRF62_8_buffer[!clk]) begin
          $fwrite(f, "Register (62,8) Value: %h\n", GRF62_8_buffer[clk]);
        end
        if (GRF62_9_buffer[clk] != GRF62_9_buffer[!clk]) begin
          $fwrite(f, "Register (62,9) Value: %h\n", GRF62_9_buffer[clk]);
        end
        if (GRF62_10_buffer[clk] != GRF62_10_buffer[!clk]) begin
          $fwrite(f, "Register (62,10) Value: %h\n", GRF62_10_buffer[clk]);
        end
        if (GRF62_11_buffer[clk] != GRF62_11_buffer[!clk]) begin
          $fwrite(f, "Register (62,11) Value: %h\n", GRF62_11_buffer[clk]);
        end
        if (GRF62_12_buffer[clk] != GRF62_12_buffer[!clk]) begin
          $fwrite(f, "Register (62,12) Value: %h\n", GRF62_12_buffer[clk]);
        end
        if (GRF62_13_buffer[clk] != GRF62_13_buffer[!clk]) begin
          $fwrite(f, "Register (62,13) Value: %h\n", GRF62_13_buffer[clk]);
        end
        if (GRF62_14_buffer[clk] != GRF62_14_buffer[!clk]) begin
          $fwrite(f, "Register (62,14) Value: %h\n", GRF62_14_buffer[clk]);
        end
        if (GRF62_15_buffer[clk] != GRF62_15_buffer[!clk]) begin
          $fwrite(f, "Register (62,15) Value: %h\n", GRF62_15_buffer[clk]);
        end
        if (GRF62_16_buffer[clk] != GRF62_16_buffer[!clk]) begin
          $fwrite(f, "Register (62,16) Value: %h\n", GRF62_16_buffer[clk]);
        end
        if (GRF62_17_buffer[clk] != GRF62_17_buffer[!clk]) begin
          $fwrite(f, "Register (62,17) Value: %h\n", GRF62_17_buffer[clk]);
        end
        if (GRF62_18_buffer[clk] != GRF62_18_buffer[!clk]) begin
          $fwrite(f, "Register (62,18) Value: %h\n", GRF62_18_buffer[clk]);
        end
        if (GRF62_19_buffer[clk] != GRF62_19_buffer[!clk]) begin
          $fwrite(f, "Register (62,19) Value: %h\n", GRF62_19_buffer[clk]);
        end
        if (GRF62_20_buffer[clk] != GRF62_20_buffer[!clk]) begin
          $fwrite(f, "Register (62,20) Value: %h\n", GRF62_20_buffer[clk]);
        end
        if (GRF62_21_buffer[clk] != GRF62_21_buffer[!clk]) begin
          $fwrite(f, "Register (62,21) Value: %h\n", GRF62_21_buffer[clk]);
        end
        if (GRF62_22_buffer[clk] != GRF62_22_buffer[!clk]) begin
          $fwrite(f, "Register (62,22) Value: %h\n", GRF62_22_buffer[clk]);
        end
        if (GRF62_23_buffer[clk] != GRF62_23_buffer[!clk]) begin
          $fwrite(f, "Register (62,23) Value: %h\n", GRF62_23_buffer[clk]);
        end
        if (GRF62_24_buffer[clk] != GRF62_24_buffer[!clk]) begin
          $fwrite(f, "Register (62,24) Value: %h\n", GRF62_24_buffer[clk]);
        end
        if (GRF62_25_buffer[clk] != GRF62_25_buffer[!clk]) begin
          $fwrite(f, "Register (62,25) Value: %h\n", GRF62_25_buffer[clk]);
        end
        if (GRF62_26_buffer[clk] != GRF62_26_buffer[!clk]) begin
          $fwrite(f, "Register (62,26) Value: %h\n", GRF62_26_buffer[clk]);
        end
        if (GRF62_27_buffer[clk] != GRF62_27_buffer[!clk]) begin
          $fwrite(f, "Register (62,27) Value: %h\n", GRF62_27_buffer[clk]);
        end
        if (GRF62_28_buffer[clk] != GRF62_28_buffer[!clk]) begin
          $fwrite(f, "Register (62,28) Value: %h\n", GRF62_28_buffer[clk]);
        end
        if (GRF62_29_buffer[clk] != GRF62_29_buffer[!clk]) begin
          $fwrite(f, "Register (62,29) Value: %h\n", GRF62_29_buffer[clk]);
        end
        if (GRF62_30_buffer[clk] != GRF62_30_buffer[!clk]) begin
          $fwrite(f, "Register (62,30) Value: %h\n", GRF62_30_buffer[clk]);
        end
        if (GRF62_31_buffer[clk] != GRF62_31_buffer[!clk]) begin
          $fwrite(f, "Register (62,31) Value: %h\n", GRF62_31_buffer[clk]);
        end
        if (GRF63_0_buffer[clk] != GRF63_0_buffer[!clk]) begin
          $fwrite(f, "Register (63,0) Value: %h\n", GRF63_0_buffer[clk]);
        end
        if (GRF63_1_buffer[clk] != GRF63_1_buffer[!clk]) begin
          $fwrite(f, "Register (63,1) Value: %h\n", GRF63_1_buffer[clk]);
        end
        if (GRF63_2_buffer[clk] != GRF63_2_buffer[!clk]) begin
          $fwrite(f, "Register (63,2) Value: %h\n", GRF63_2_buffer[clk]);
        end
        if (GRF63_3_buffer[clk] != GRF63_3_buffer[!clk]) begin
          $fwrite(f, "Register (63,3) Value: %h\n", GRF63_3_buffer[clk]);
        end
        if (GRF63_4_buffer[clk] != GRF63_4_buffer[!clk]) begin
          $fwrite(f, "Register (63,4) Value: %h\n", GRF63_4_buffer[clk]);
        end
        if (GRF63_5_buffer[clk] != GRF63_5_buffer[!clk]) begin
          $fwrite(f, "Register (63,5) Value: %h\n", GRF63_5_buffer[clk]);
        end
        if (GRF63_6_buffer[clk] != GRF63_6_buffer[!clk]) begin
          $fwrite(f, "Register (63,6) Value: %h\n", GRF63_6_buffer[clk]);
        end
        if (GRF63_7_buffer[clk] != GRF63_7_buffer[!clk]) begin
          $fwrite(f, "Register (63,7) Value: %h\n", GRF63_7_buffer[clk]);
        end
        if (GRF63_8_buffer[clk] != GRF63_8_buffer[!clk]) begin
          $fwrite(f, "Register (63,8) Value: %h\n", GRF63_8_buffer[clk]);
        end
        if (GRF63_9_buffer[clk] != GRF63_9_buffer[!clk]) begin
          $fwrite(f, "Register (63,9) Value: %h\n", GRF63_9_buffer[clk]);
        end
        if (GRF63_10_buffer[clk] != GRF63_10_buffer[!clk]) begin
          $fwrite(f, "Register (63,10) Value: %h\n", GRF63_10_buffer[clk]);
        end
        if (GRF63_11_buffer[clk] != GRF63_11_buffer[!clk]) begin
          $fwrite(f, "Register (63,11) Value: %h\n", GRF63_11_buffer[clk]);
        end
        if (GRF63_12_buffer[clk] != GRF63_12_buffer[!clk]) begin
          $fwrite(f, "Register (63,12) Value: %h\n", GRF63_12_buffer[clk]);
        end
        if (GRF63_13_buffer[clk] != GRF63_13_buffer[!clk]) begin
          $fwrite(f, "Register (63,13) Value: %h\n", GRF63_13_buffer[clk]);
        end
        if (GRF63_14_buffer[clk] != GRF63_14_buffer[!clk]) begin
          $fwrite(f, "Register (63,14) Value: %h\n", GRF63_14_buffer[clk]);
        end
        if (GRF63_15_buffer[clk] != GRF63_15_buffer[!clk]) begin
          $fwrite(f, "Register (63,15) Value: %h\n", GRF63_15_buffer[clk]);
        end
        if (GRF63_16_buffer[clk] != GRF63_16_buffer[!clk]) begin
          $fwrite(f, "Register (63,16) Value: %h\n", GRF63_16_buffer[clk]);
        end
        if (GRF63_17_buffer[clk] != GRF63_17_buffer[!clk]) begin
          $fwrite(f, "Register (63,17) Value: %h\n", GRF63_17_buffer[clk]);
        end
        if (GRF63_18_buffer[clk] != GRF63_18_buffer[!clk]) begin
          $fwrite(f, "Register (63,18) Value: %h\n", GRF63_18_buffer[clk]);
        end
        if (GRF63_19_buffer[clk] != GRF63_19_buffer[!clk]) begin
          $fwrite(f, "Register (63,19) Value: %h\n", GRF63_19_buffer[clk]);
        end
        if (GRF63_20_buffer[clk] != GRF63_20_buffer[!clk]) begin
          $fwrite(f, "Register (63,20) Value: %h\n", GRF63_20_buffer[clk]);
        end
        if (GRF63_21_buffer[clk] != GRF63_21_buffer[!clk]) begin
          $fwrite(f, "Register (63,21) Value: %h\n", GRF63_21_buffer[clk]);
        end
        if (GRF63_22_buffer[clk] != GRF63_22_buffer[!clk]) begin
          $fwrite(f, "Register (63,22) Value: %h\n", GRF63_22_buffer[clk]);
        end
        if (GRF63_23_buffer[clk] != GRF63_23_buffer[!clk]) begin
          $fwrite(f, "Register (63,23) Value: %h\n", GRF63_23_buffer[clk]);
        end
        if (GRF63_24_buffer[clk] != GRF63_24_buffer[!clk]) begin
          $fwrite(f, "Register (63,24) Value: %h\n", GRF63_24_buffer[clk]);
        end
        if (GRF63_25_buffer[clk] != GRF63_25_buffer[!clk]) begin
          $fwrite(f, "Register (63,25) Value: %h\n", GRF63_25_buffer[clk]);
        end
        if (GRF63_26_buffer[clk] != GRF63_26_buffer[!clk]) begin
          $fwrite(f, "Register (63,26) Value: %h\n", GRF63_26_buffer[clk]);
        end
        if (GRF63_27_buffer[clk] != GRF63_27_buffer[!clk]) begin
          $fwrite(f, "Register (63,27) Value: %h\n", GRF63_27_buffer[clk]);
        end
        if (GRF63_28_buffer[clk] != GRF63_28_buffer[!clk]) begin
          $fwrite(f, "Register (63,28) Value: %h\n", GRF63_28_buffer[clk]);
        end
        if (GRF63_29_buffer[clk] != GRF63_29_buffer[!clk]) begin
          $fwrite(f, "Register (63,29) Value: %h\n", GRF63_29_buffer[clk]);
        end
        if (GRF63_30_buffer[clk] != GRF63_30_buffer[!clk]) begin
          $fwrite(f, "Register (63,30) Value: %h\n", GRF63_30_buffer[clk]);
        end
        if (GRF63_31_buffer[clk] != GRF63_31_buffer[!clk]) begin
          $fwrite(f, "Register (63,31) Value: %h\n", GRF63_31_buffer[clk]);
        end

        $fwrite(f, " \n=====================================================\n\n\n\n\n");
      end
    end
    $fclose(f);
  end 

endmodule









